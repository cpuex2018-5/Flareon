`timescale 1ns / 1ps

//とりあえず組み合わせ回路で実現しようか
//s<0に対しては出力てきとう

//以下、すごく注意なのだが、
//まずは入力xに対してx^(-1/2)を求め、これにxをかけてsqrt(x)を求めることにしているよ

module fsqrt(
  input clk,
  input [31:0] x,
  output [31:0] y);
  
  wire sx;
  wire [7:0] ex;
  wire [22:0] mx;
  
  assign {sx,ex,mx}=x;
  
  //25bit_verに対応させた
  wire [25:0] three;
  wire [25:0] cube;

  logic [25:0] three_reg;
  logic [25:0] cube_reg;
  
  //テーブルをもとに作成
  assign three = 
  (x[23:13] == 0) ? 26'b10000111101110110011101100 :
  (x[23:13] == 1) ? 26'b10000111101010100100100100 :
  (x[23:13] == 2) ? 26'b10000111100110010101110100 :
  (x[23:13] == 3) ? 26'b10000111100010000111100000 :
  (x[23:13] == 4) ? 26'b10000111011101111001100000 :
  (x[23:13] == 5) ? 26'b10000111011001101100000000 :
  (x[23:13] == 6) ? 26'b10000111010101011110110100 :
  (x[23:13] == 7) ? 26'b10000111010001010010000100 :
  (x[23:13] == 8) ? 26'b10000111001101000101101000 :
  (x[23:13] == 9) ? 26'b10000111001000111001101100 :
  (x[23:13] == 10) ? 26'b10000111000100101110000100 :
  (x[23:13] == 11) ? 26'b10000111000000100010111000 :
  (x[23:13] == 12) ? 26'b10000110111100011000000100 :
  (x[23:13] == 13) ? 26'b10000110111000001101101000 :
  (x[23:13] == 14) ? 26'b10000110110100000011100100 :
  (x[23:13] == 15) ? 26'b10000110101111111001111000 :
  (x[23:13] == 16) ? 26'b10000110101011110000101000 :
  (x[23:13] == 17) ? 26'b10000110100111100111101100 :
  (x[23:13] == 18) ? 26'b10000110100011011111001000 :
  (x[23:13] == 19) ? 26'b10000110011111010111000000 :
  (x[23:13] == 20) ? 26'b10000110011011001111010000 :
  (x[23:13] == 21) ? 26'b10000110010111000111111000 :
  (x[23:13] == 22) ? 26'b10000110010011000000111000 :
  (x[23:13] == 23) ? 26'b10000110001110111010010000 :
  (x[23:13] == 24) ? 26'b10000110001010110100000000 :
  (x[23:13] == 25) ? 26'b10000110000110101110001000 :
  (x[23:13] == 26) ? 26'b10000110000010101000100100 :
  (x[23:13] == 27) ? 26'b10000101111110100011100000 :
  (x[23:13] == 28) ? 26'b10000101111010011110110000 :
  (x[23:13] == 29) ? 26'b10000101110110011010010100 :
  (x[23:13] == 30) ? 26'b10000101110010010110010100 :
  (x[23:13] == 31) ? 26'b10000101101110010010101000 :
  (x[23:13] == 32) ? 26'b10000101101010001111011000 :
  (x[23:13] == 33) ? 26'b10000101100110001100100000 :
  (x[23:13] == 34) ? 26'b10000101100010001001111000 :
  (x[23:13] == 35) ? 26'b10000101011110000111110000 :
  (x[23:13] == 36) ? 26'b10000101011010000101111000 :
  (x[23:13] == 37) ? 26'b10000101010110000100100000 :
  (x[23:13] == 38) ? 26'b10000101010010000011011000 :
  (x[23:13] == 39) ? 26'b10000101001110000010101000 :
  (x[23:13] == 40) ? 26'b10000101001010000010010000 :
  (x[23:13] == 41) ? 26'b10000101000110000010010000 :
  (x[23:13] == 42) ? 26'b10000101000010000010101000 :
  (x[23:13] == 43) ? 26'b10000100111110000011011000 :
  (x[23:13] == 44) ? 26'b10000100111010000100011100 :
  (x[23:13] == 45) ? 26'b10000100110110000101111000 :
  (x[23:13] == 46) ? 26'b10000100110010000111101000 :
  (x[23:13] == 47) ? 26'b10000100101110001001110100 :
  (x[23:13] == 48) ? 26'b10000100101010001100010100 :
  (x[23:13] == 49) ? 26'b10000100100110001111001000 :
  (x[23:13] == 50) ? 26'b10000100100010010010011000 :
  (x[23:13] == 51) ? 26'b10000100011110010101111100 :
  (x[23:13] == 52) ? 26'b10000100011010011001111000 :
  (x[23:13] == 53) ? 26'b10000100010110011110001000 :
  (x[23:13] == 54) ? 26'b10000100010010100010110000 :
  (x[23:13] == 55) ? 26'b10000100001110100111110000 :
  (x[23:13] == 56) ? 26'b10000100001010101101000000 :
  (x[23:13] == 57) ? 26'b10000100000110110010101100 :
  (x[23:13] == 58) ? 26'b10000100000010111000101100 :
  (x[23:13] == 59) ? 26'b10000011111110111111000000 :
  (x[23:13] == 60) ? 26'b10000011111011000101110000 :
  (x[23:13] == 61) ? 26'b10000011110111001100110100 :
  (x[23:13] == 62) ? 26'b10000011110011010100001100 :
  (x[23:13] == 63) ? 26'b10000011101111011011111100 :
  (x[23:13] == 64) ? 26'b10000011101011100100000000 :
  (x[23:13] == 65) ? 26'b10000011100111101100011000 :
  (x[23:13] == 66) ? 26'b10000011100011110101001000 :
  (x[23:13] == 67) ? 26'b10000011011111111110010000 :
  (x[23:13] == 68) ? 26'b10000011011100000111101100 :
  (x[23:13] == 69) ? 26'b10000011011000010001011100 :
  (x[23:13] == 70) ? 26'b10000011010100011011100100 :
  (x[23:13] == 71) ? 26'b10000011010000100110000000 :
  (x[23:13] == 72) ? 26'b10000011001100110000110100 :
  (x[23:13] == 73) ? 26'b10000011001000111011111000 :
  (x[23:13] == 74) ? 26'b10000011000101000111011000 :
  (x[23:13] == 75) ? 26'b10000011000001010011001100 :
  (x[23:13] == 76) ? 26'b10000010111101011111010000 :
  (x[23:13] == 77) ? 26'b10000010111001101011110000 :
  (x[23:13] == 78) ? 26'b10000010110101111000100000 :
  (x[23:13] == 79) ? 26'b10000010110010000101101000 :
  (x[23:13] == 80) ? 26'b10000010101110010011000100 :
  (x[23:13] == 81) ? 26'b10000010101010100000111000 :
  (x[23:13] == 82) ? 26'b10000010100110101110111100 :
  (x[23:13] == 83) ? 26'b10000010100010111101011000 :
  (x[23:13] == 84) ? 26'b10000010011111001100001000 :
  (x[23:13] == 85) ? 26'b10000010011011011011010000 :
  (x[23:13] == 86) ? 26'b10000010010111101010101000 :
  (x[23:13] == 87) ? 26'b10000010010011111010010100 :
  (x[23:13] == 88) ? 26'b10000010010000001010011100 :
  (x[23:13] == 89) ? 26'b10000010001100011010110100 :
  (x[23:13] == 90) ? 26'b10000010001000101011100000 :
  (x[23:13] == 91) ? 26'b10000010000100111100100000 :
  (x[23:13] == 92) ? 26'b10000010000001001101111000 :
  (x[23:13] == 93) ? 26'b10000001111101011111100000 :
  (x[23:13] == 94) ? 26'b10000001111001110001100000 :
  (x[23:13] == 95) ? 26'b10000001110110000011110100 :
  (x[23:13] == 96) ? 26'b10000001110010010110011100 :
  (x[23:13] == 97) ? 26'b10000001101110101001011000 :
  (x[23:13] == 98) ? 26'b10000001101010111100101000 :
  (x[23:13] == 99) ? 26'b10000001100111010000010000 :
  (x[23:13] == 100) ? 26'b10000001100011100100001000 :
  (x[23:13] == 101) ? 26'b10000001011111111000010000 :
  (x[23:13] == 102) ? 26'b10000001011100001100110100 :
  (x[23:13] == 103) ? 26'b10000001011000100001101000 :
  (x[23:13] == 104) ? 26'b10000001010100110110110000 :
  (x[23:13] == 105) ? 26'b10000001010001001100010000 :
  (x[23:13] == 106) ? 26'b10000001001101100010000000 :
  (x[23:13] == 107) ? 26'b10000001001001111000001000 :
  (x[23:13] == 108) ? 26'b10000001000110001110100000 :
  (x[23:13] == 109) ? 26'b10000001000010100101001100 :
  (x[23:13] == 110) ? 26'b10000000111110111100001100 :
  (x[23:13] == 111) ? 26'b10000000111011010011100000 :
  (x[23:13] == 112) ? 26'b10000000110111101011001000 :
  (x[23:13] == 113) ? 26'b10000000110100000011000100 :
  (x[23:13] == 114) ? 26'b10000000110000011011010000 :
  (x[23:13] == 115) ? 26'b10000000101100110011110000 :
  (x[23:13] == 116) ? 26'b10000000101001001100101000 :
  (x[23:13] == 117) ? 26'b10000000100101100101110000 :
  (x[23:13] == 118) ? 26'b10000000100001111111010000 :
  (x[23:13] == 119) ? 26'b10000000011110011001000000 :
  (x[23:13] == 120) ? 26'b10000000011010110011000000 :
  (x[23:13] == 121) ? 26'b10000000010111001101011000 :
  (x[23:13] == 122) ? 26'b10000000010011101000000100 :
  (x[23:13] == 123) ? 26'b10000000010000000011000000 :
  (x[23:13] == 124) ? 26'b10000000001100011110010000 :
  (x[23:13] == 125) ? 26'b10000000001000111001110100 :
  (x[23:13] == 126) ? 26'b10000000000101010101101100 :
  (x[23:13] == 127) ? 26'b10000000000001110001110100 :
  (x[23:13] == 128) ? 26'b01111111111110001110010000 :
  (x[23:13] == 129) ? 26'b01111111111010101011000000 :
  (x[23:13] == 130) ? 26'b01111111110111001000000010 :
  (x[23:13] == 131) ? 26'b01111111110011100101010110 :
  (x[23:13] == 132) ? 26'b01111111110000000011000000 :
  (x[23:13] == 133) ? 26'b01111111101100100000111010 :
  (x[23:13] == 134) ? 26'b01111111101000111111001000 :
  (x[23:13] == 135) ? 26'b01111111100101011101101000 :
  (x[23:13] == 136) ? 26'b01111111100001111100011010 :
  (x[23:13] == 137) ? 26'b01111111011110011011100000 :
  (x[23:13] == 138) ? 26'b01111111011010111010111000 :
  (x[23:13] == 139) ? 26'b01111111010111011010100010 :
  (x[23:13] == 140) ? 26'b01111111010011111010100000 :
  (x[23:13] == 141) ? 26'b01111111010000011010110000 :
  (x[23:13] == 142) ? 26'b01111111001100111011010010 :
  (x[23:13] == 143) ? 26'b01111111001001011100001000 :
  (x[23:13] == 144) ? 26'b01111111000101111101001100 :
  (x[23:13] == 145) ? 26'b01111111000010011110100100 :
  (x[23:13] == 146) ? 26'b01111110111111000000010000 :
  (x[23:13] == 147) ? 26'b01111110111011100010010000 :
  (x[23:13] == 148) ? 26'b01111110111000000100011110 :
  (x[23:13] == 149) ? 26'b01111110110100100111000000 :
  (x[23:13] == 150) ? 26'b01111110110001001001110010 :
  (x[23:13] == 151) ? 26'b01111110101101101100111010 :
  (x[23:13] == 152) ? 26'b01111110101010010000010000 :
  (x[23:13] == 153) ? 26'b01111110100110110011111010 :
  (x[23:13] == 154) ? 26'b01111110100011010111111000 :
  (x[23:13] == 155) ? 26'b01111110011111111100000100 :
  (x[23:13] == 156) ? 26'b01111110011100100000100100 :
  (x[23:13] == 157) ? 26'b01111110011001000101010100 :
  (x[23:13] == 158) ? 26'b01111110010101101010011100 :
  (x[23:13] == 159) ? 26'b01111110010010001111110000 :
  (x[23:13] == 160) ? 26'b01111110001110110101010100 :
  (x[23:13] == 161) ? 26'b01111110001011011011001100 :
  (x[23:13] == 162) ? 26'b01111110001000000001011000 :
  (x[23:13] == 163) ? 26'b01111110000100100111110100 :
  (x[23:13] == 164) ? 26'b01111110000001001110100000 :
  (x[23:13] == 165) ? 26'b01111101111101110101100000 :
  (x[23:13] == 166) ? 26'b01111101111010011100110010 :
  (x[23:13] == 167) ? 26'b01111101110111000100010100 :
  (x[23:13] == 168) ? 26'b01111101110011101100000100 :
  (x[23:13] == 169) ? 26'b01111101110000010100001100 :
  (x[23:13] == 170) ? 26'b01111101101100111100100000 :
  (x[23:13] == 171) ? 26'b01111101101001100101001000 :
  (x[23:13] == 172) ? 26'b01111101100110001110000000 :
  (x[23:13] == 173) ? 26'b01111101100010110111001100 :
  (x[23:13] == 174) ? 26'b01111101011111100000100100 :
  (x[23:13] == 175) ? 26'b01111101011100001010010000 :
  (x[23:13] == 176) ? 26'b01111101011000110100010000 :
  (x[23:13] == 177) ? 26'b01111101010101011110100000 :
  (x[23:13] == 178) ? 26'b01111101010010001000111110 :
  (x[23:13] == 179) ? 26'b01111101001110110011110000 :
  (x[23:13] == 180) ? 26'b01111101001011011110110000 :
  (x[23:13] == 181) ? 26'b01111101001000001010000100 :
  (x[23:13] == 182) ? 26'b01111101000100110101100100 :
  (x[23:13] == 183) ? 26'b01111101000001100001011100 :
  (x[23:13] == 184) ? 26'b01111100111110001101100000 :
  (x[23:13] == 185) ? 26'b01111100111010111001111000 :
  (x[23:13] == 186) ? 26'b01111100110111100110011100 :
  (x[23:13] == 187) ? 26'b01111100110100010011010100 :
  (x[23:13] == 188) ? 26'b01111100110001000000011100 :
  (x[23:13] == 189) ? 26'b01111100101101101101110100 :
  (x[23:13] == 190) ? 26'b01111100101010011011100000 :
  (x[23:13] == 191) ? 26'b01111100100111001001011010 :
  (x[23:13] == 192) ? 26'b01111100100011110111100110 :
  (x[23:13] == 193) ? 26'b01111100100000100110000000 :
  (x[23:13] == 194) ? 26'b01111100011101010100101110 :
  (x[23:13] == 195) ? 26'b01111100011010000011101010 :
  (x[23:13] == 196) ? 26'b01111100010110110010110100 :
  (x[23:13] == 197) ? 26'b01111100010011100010010100 :
  (x[23:13] == 198) ? 26'b01111100010000010010000000 :
  (x[23:13] == 199) ? 26'b01111100001101000010000000 :
  (x[23:13] == 200) ? 26'b01111100001001110010010000 :
  (x[23:13] == 201) ? 26'b01111100000110100010101100 :
  (x[23:13] == 202) ? 26'b01111100000011010011011100 :
  (x[23:13] == 203) ? 26'b01111100000000000100011000 :
  (x[23:13] == 204) ? 26'b01111011111100110101101100 :
  (x[23:13] == 205) ? 26'b01111011111001100111001000 :
  (x[23:13] == 206) ? 26'b01111011110110011000111000 :
  (x[23:13] == 207) ? 26'b01111011110011001010111000 :
  (x[23:13] == 208) ? 26'b01111011101111111101001000 :
  (x[23:13] == 209) ? 26'b01111011101100101111101000 :
  (x[23:13] == 210) ? 26'b01111011101001100010011000 :
  (x[23:13] == 211) ? 26'b01111011100110010101010110 :
  (x[23:13] == 212) ? 26'b01111011100011001000100110 :
  (x[23:13] == 213) ? 26'b01111011011111111100000100 :
  (x[23:13] == 214) ? 26'b01111011011100101111110110 :
  (x[23:13] == 215) ? 26'b01111011011001100011110110 :
  (x[23:13] == 216) ? 26'b01111011010110011000000010 :
  (x[23:13] == 217) ? 26'b01111011010011001100100100 :
  (x[23:13] == 218) ? 26'b01111011010000000001010000 :
  (x[23:13] == 219) ? 26'b01111011001100110110010000 :
  (x[23:13] == 220) ? 26'b01111011001001101011011100 :
  (x[23:13] == 221) ? 26'b01111011000110100000111010 :
  (x[23:13] == 222) ? 26'b01111011000011010110100110 :
  (x[23:13] == 223) ? 26'b01111011000000001100100100 :
  (x[23:13] == 224) ? 26'b01111010111101000010101110 :
  (x[23:13] == 225) ? 26'b01111010111001111001001010 :
  (x[23:13] == 226) ? 26'b01111010110110101111110100 :
  (x[23:13] == 227) ? 26'b01111010110011100110110010 :
  (x[23:13] == 228) ? 26'b01111010110000011101111100 :
  (x[23:13] == 229) ? 26'b01111010101101010101010100 :
  (x[23:13] == 230) ? 26'b01111010101010001100111100 :
  (x[23:13] == 231) ? 26'b01111010100111000100110110 :
  (x[23:13] == 232) ? 26'b01111010100011111100111100 :
  (x[23:13] == 233) ? 26'b01111010100000110101010010 :
  (x[23:13] == 234) ? 26'b01111010011101101101111000 :
  (x[23:13] == 235) ? 26'b01111010011010100110101100 :
  (x[23:13] == 236) ? 26'b01111010010111011111110000 :
  (x[23:13] == 237) ? 26'b01111010010100011001000100 :
  (x[23:13] == 238) ? 26'b01111010010001010010100110 :
  (x[23:13] == 239) ? 26'b01111010001110001100011010 :
  (x[23:13] == 240) ? 26'b01111010001011000110011010 :
  (x[23:13] == 241) ? 26'b01111010001000000000101000 :
  (x[23:13] == 242) ? 26'b01111010000100111011001000 :
  (x[23:13] == 243) ? 26'b01111010000001110101110100 :
  (x[23:13] == 244) ? 26'b01111001111110110000110100 :
  (x[23:13] == 245) ? 26'b01111001111011101011111110 :
  (x[23:13] == 246) ? 26'b01111001111000100111011000 :
  (x[23:13] == 247) ? 26'b01111001110101100011000000 :
  (x[23:13] == 248) ? 26'b01111001110010011110111000 :
  (x[23:13] == 249) ? 26'b01111001101111011011000000 :
  (x[23:13] == 250) ? 26'b01111001101100010111010110 :
  (x[23:13] == 251) ? 26'b01111001101001010011111000 :
  (x[23:13] == 252) ? 26'b01111001100110010000101100 :
  (x[23:13] == 253) ? 26'b01111001100011001101101100 :
  (x[23:13] == 254) ? 26'b01111001100000001010111110 :
  (x[23:13] == 255) ? 26'b01111001011101001000011100 :
  (x[23:13] == 256) ? 26'b01111001011010000110001000 :
  (x[23:13] == 257) ? 26'b01111001010111000100000100 :
  (x[23:13] == 258) ? 26'b01111001010100000010010000 :
  (x[23:13] == 259) ? 26'b01111001010001000000101010 :
  (x[23:13] == 260) ? 26'b01111001001101111111010000 :
  (x[23:13] == 261) ? 26'b01111001001010111110001000 :
  (x[23:13] == 262) ? 26'b01111001000111111101001100 :
  (x[23:13] == 263) ? 26'b01111001000100111100100000 :
  (x[23:13] == 264) ? 26'b01111001000001111011111110 :
  (x[23:13] == 265) ? 26'b01111000111110111011110000 :
  (x[23:13] == 266) ? 26'b01111000111011111011101100 :
  (x[23:13] == 267) ? 26'b01111000111000111011111000 :
  (x[23:13] == 268) ? 26'b01111000110101111100010100 :
  (x[23:13] == 269) ? 26'b01111000110010111100111010 :
  (x[23:13] == 270) ? 26'b01111000101111111101110000 :
  (x[23:13] == 271) ? 26'b01111000101100111110110100 :
  (x[23:13] == 272) ? 26'b01111000101010000000001000 :
  (x[23:13] == 273) ? 26'b01111000100111000001101000 :
  (x[23:13] == 274) ? 26'b01111000100100000011011000 :
  (x[23:13] == 275) ? 26'b01111000100001000101010110 :
  (x[23:13] == 276) ? 26'b01111000011110000111100100 :
  (x[23:13] == 277) ? 26'b01111000011011001001111100 :
  (x[23:13] == 278) ? 26'b01111000011000001100100000 :
  (x[23:13] == 279) ? 26'b01111000010101001111011000 :
  (x[23:13] == 280) ? 26'b01111000010010010010011100 :
  (x[23:13] == 281) ? 26'b01111000001111010101101100 :
  (x[23:13] == 282) ? 26'b01111000001100011001001100 :
  (x[23:13] == 283) ? 26'b01111000001001011100111000 :
  (x[23:13] == 284) ? 26'b01111000000110100000110000 :
  (x[23:13] == 285) ? 26'b01111000000011100100111000 :
  (x[23:13] == 286) ? 26'b01111000000000101001010000 :
  (x[23:13] == 287) ? 26'b01110111111101101101110100 :
  (x[23:13] == 288) ? 26'b01110111111010110010100100 :
  (x[23:13] == 289) ? 26'b01110111110111110111100110 :
  (x[23:13] == 290) ? 26'b01110111110100111100110100 :
  (x[23:13] == 291) ? 26'b01110111110010000010001100 :
  (x[23:13] == 292) ? 26'b01110111101111000111110100 :
  (x[23:13] == 293) ? 26'b01110111101100001101101100 :
  (x[23:13] == 294) ? 26'b01110111101001010011101110 :
  (x[23:13] == 295) ? 26'b01110111100110011001111100 :
  (x[23:13] == 296) ? 26'b01110111100011100000011110 :
  (x[23:13] == 297) ? 26'b01110111100000100111001000 :
  (x[23:13] == 298) ? 26'b01110111011101101110000000 :
  (x[23:13] == 299) ? 26'b01110111011010110101001000 :
  (x[23:13] == 300) ? 26'b01110111010111111100011100 :
  (x[23:13] == 301) ? 26'b01110111010101000011111100 :
  (x[23:13] == 302) ? 26'b01110111010010001011101100 :
  (x[23:13] == 303) ? 26'b01110111001111010011101010 :
  (x[23:13] == 304) ? 26'b01110111001100011011110000 :
  (x[23:13] == 305) ? 26'b01110111001001100100001010 :
  (x[23:13] == 306) ? 26'b01110111000110101100101100 :
  (x[23:13] == 307) ? 26'b01110111000011110101011100 :
  (x[23:13] == 308) ? 26'b01110111000000111110011100 :
  (x[23:13] == 309) ? 26'b01110110111110000111101000 :
  (x[23:13] == 310) ? 26'b01110110111011010001000000 :
  (x[23:13] == 311) ? 26'b01110110111000011010101000 :
  (x[23:13] == 312) ? 26'b01110110110101100100011100 :
  (x[23:13] == 313) ? 26'b01110110110010101110011010 :
  (x[23:13] == 314) ? 26'b01110110101111111000101000 :
  (x[23:13] == 315) ? 26'b01110110101101000011000010 :
  (x[23:13] == 316) ? 26'b01110110101010001101101000 :
  (x[23:13] == 317) ? 26'b01110110100111011000011100 :
  (x[23:13] == 318) ? 26'b01110110100100100011011110 :
  (x[23:13] == 319) ? 26'b01110110100001101110101100 :
  (x[23:13] == 320) ? 26'b01110110011110111010001000 :
  (x[23:13] == 321) ? 26'b01110110011100000101110000 :
  (x[23:13] == 322) ? 26'b01110110011001010001100100 :
  (x[23:13] == 323) ? 26'b01110110010110011101100110 :
  (x[23:13] == 324) ? 26'b01110110010011101001110010 :
  (x[23:13] == 325) ? 26'b01110110010000110110001100 :
  (x[23:13] == 326) ? 26'b01110110001110000010111000 :
  (x[23:13] == 327) ? 26'b01110110001011001111101010 :
  (x[23:13] == 328) ? 26'b01110110001000011100101100 :
  (x[23:13] == 329) ? 26'b01110110000101101001111010 :
  (x[23:13] == 330) ? 26'b01110110000010110111010100 :
  (x[23:13] == 331) ? 26'b01110110000000000100111100 :
  (x[23:13] == 332) ? 26'b01110101111101010010110000 :
  (x[23:13] == 333) ? 26'b01110101111010100000110000 :
  (x[23:13] == 334) ? 26'b01110101110111101110111100 :
  (x[23:13] == 335) ? 26'b01110101110100111101011000 :
  (x[23:13] == 336) ? 26'b01110101110010001011111110 :
  (x[23:13] == 337) ? 26'b01110101101111011010110010 :
  (x[23:13] == 338) ? 26'b01110101101100101001110000 :
  (x[23:13] == 339) ? 26'b01110101101001111000111100 :
  (x[23:13] == 340) ? 26'b01110101100111001000010100 :
  (x[23:13] == 341) ? 26'b01110101100100010111111010 :
  (x[23:13] == 342) ? 26'b01110101100001100111101010 :
  (x[23:13] == 343) ? 26'b01110101011110110111100110 :
  (x[23:13] == 344) ? 26'b01110101011100000111110000 :
  (x[23:13] == 345) ? 26'b01110101011001011000001000 :
  (x[23:13] == 346) ? 26'b01110101010110101000101000 :
  (x[23:13] == 347) ? 26'b01110101010011111001011000 :
  (x[23:13] == 348) ? 26'b01110101010001001010010010 :
  (x[23:13] == 349) ? 26'b01110101001110011011011000 :
  (x[23:13] == 350) ? 26'b01110101001011101100110000 :
  (x[23:13] == 351) ? 26'b01110101001000111110001110 :
  (x[23:13] == 352) ? 26'b01110101000110001111111000 :
  (x[23:13] == 353) ? 26'b01110101000011100001110000 :
  (x[23:13] == 354) ? 26'b01110101000000110011110110 :
  (x[23:13] == 355) ? 26'b01110100111110000110000100 :
  (x[23:13] == 356) ? 26'b01110100111011011000100000 :
  (x[23:13] == 357) ? 26'b01110100111000101011001010 :
  (x[23:13] == 358) ? 26'b01110100110101111101111100 :
  (x[23:13] == 359) ? 26'b01110100110011010001000000 :
  (x[23:13] == 360) ? 26'b01110100110000100100001010 :
  (x[23:13] == 361) ? 26'b01110100101101110111100100 :
  (x[23:13] == 362) ? 26'b01110100101011001011001000 :
  (x[23:13] == 363) ? 26'b01110100101000011110110110 :
  (x[23:13] == 364) ? 26'b01110100100101110010110100 :
  (x[23:13] == 365) ? 26'b01110100100011000110111100 :
  (x[23:13] == 366) ? 26'b01110100100000011011001110 :
  (x[23:13] == 367) ? 26'b01110100011101101111110000 :
  (x[23:13] == 368) ? 26'b01110100011011000100011100 :
  (x[23:13] == 369) ? 26'b01110100011000011001010010 :
  (x[23:13] == 370) ? 26'b01110100010101101110010100 :
  (x[23:13] == 371) ? 26'b01110100010011000011100100 :
  (x[23:13] == 372) ? 26'b01110100010000011001000000 :
  (x[23:13] == 373) ? 26'b01110100001101101110100110 :
  (x[23:13] == 374) ? 26'b01110100001011000100010110 :
  (x[23:13] == 375) ? 26'b01110100001000011010010100 :
  (x[23:13] == 376) ? 26'b01110100000101110000011100 :
  (x[23:13] == 377) ? 26'b01110100000011000110110100 :
  (x[23:13] == 378) ? 26'b01110100000000011101010100 :
  (x[23:13] == 379) ? 26'b01110011111101110100000000 :
  (x[23:13] == 380) ? 26'b01110011111011001010111000 :
  (x[23:13] == 381) ? 26'b01110011111000100001111100 :
  (x[23:13] == 382) ? 26'b01110011110101111001001000 :
  (x[23:13] == 383) ? 26'b01110011110011010000100100 :
  (x[23:13] == 384) ? 26'b01110011110000101000001010 :
  (x[23:13] == 385) ? 26'b01110011101101111111111100 :
  (x[23:13] == 386) ? 26'b01110011101011010111111000 :
  (x[23:13] == 387) ? 26'b01110011101000110000000000 :
  (x[23:13] == 388) ? 26'b01110011100110001000010100 :
  (x[23:13] == 389) ? 26'b01110011100011100000110100 :
  (x[23:13] == 390) ? 26'b01110011100000111001011110 :
  (x[23:13] == 391) ? 26'b01110011011110010010010100 :
  (x[23:13] == 392) ? 26'b01110011011011101011010110 :
  (x[23:13] == 393) ? 26'b01110011011001000100100000 :
  (x[23:13] == 394) ? 26'b01110011010110011101111000 :
  (x[23:13] == 395) ? 26'b01110011010011110111011100 :
  (x[23:13] == 396) ? 26'b01110011010001010001001010 :
  (x[23:13] == 397) ? 26'b01110011001110101011000010 :
  (x[23:13] == 398) ? 26'b01110011001100000101001000 :
  (x[23:13] == 399) ? 26'b01110011001001011111011000 :
  (x[23:13] == 400) ? 26'b01110011000110111001110010 :
  (x[23:13] == 401) ? 26'b01110011000100010100011010 :
  (x[23:13] == 402) ? 26'b01110011000001101111001100 :
  (x[23:13] == 403) ? 26'b01110010111111001010001000 :
  (x[23:13] == 404) ? 26'b01110010111100100101001110 :
  (x[23:13] == 405) ? 26'b01110010111010000000100000 :
  (x[23:13] == 406) ? 26'b01110010110111011011111110 :
  (x[23:13] == 407) ? 26'b01110010110100110111101000 :
  (x[23:13] == 408) ? 26'b01110010110010010011011100 :
  (x[23:13] == 409) ? 26'b01110010101111101111011010 :
  (x[23:13] == 410) ? 26'b01110010101101001011100100 :
  (x[23:13] == 411) ? 26'b01110010101010100111111000 :
  (x[23:13] == 412) ? 26'b01110010101000000100011000 :
  (x[23:13] == 413) ? 26'b01110010100101100001000010 :
  (x[23:13] == 414) ? 26'b01110010100010111101111000 :
  (x[23:13] == 415) ? 26'b01110010100000011010111000 :
  (x[23:13] == 416) ? 26'b01110010011101111000000010 :
  (x[23:13] == 417) ? 26'b01110010011011010101011000 :
  (x[23:13] == 418) ? 26'b01110010011000110010111010 :
  (x[23:13] == 419) ? 26'b01110010010110010000100100 :
  (x[23:13] == 420) ? 26'b01110010010011101110011100 :
  (x[23:13] == 421) ? 26'b01110010010001001100011100 :
  (x[23:13] == 422) ? 26'b01110010001110101010101000 :
  (x[23:13] == 423) ? 26'b01110010001100001001000000 :
  (x[23:13] == 424) ? 26'b01110010001001100111100000 :
  (x[23:13] == 425) ? 26'b01110010000111000110001110 :
  (x[23:13] == 426) ? 26'b01110010000100100101000100 :
  (x[23:13] == 427) ? 26'b01110010000010000100000110 :
  (x[23:13] == 428) ? 26'b01110001111111100011010000 :
  (x[23:13] == 429) ? 26'b01110001111101000010101000 :
  (x[23:13] == 430) ? 26'b01110001111010100010001100 :
  (x[23:13] == 431) ? 26'b01110001111000000001111000 :
  (x[23:13] == 432) ? 26'b01110001110101100001101100 :
  (x[23:13] == 433) ? 26'b01110001110011000001101100 :
  (x[23:13] == 434) ? 26'b01110001110000100001111010 :
  (x[23:13] == 435) ? 26'b01110001101110000010010000 :
  (x[23:13] == 436) ? 26'b01110001101011100010110000 :
  (x[23:13] == 437) ? 26'b01110001101001000011011010 :
  (x[23:13] == 438) ? 26'b01110001100110100100010000 :
  (x[23:13] == 439) ? 26'b01110001100100000101010000 :
  (x[23:13] == 440) ? 26'b01110001100001100110011010 :
  (x[23:13] == 441) ? 26'b01110001011111000111110000 :
  (x[23:13] == 442) ? 26'b01110001011100101001001100 :
  (x[23:13] == 443) ? 26'b01110001011010001010111000 :
  (x[23:13] == 444) ? 26'b01110001010111101100101100 :
  (x[23:13] == 445) ? 26'b01110001010101001110101000 :
  (x[23:13] == 446) ? 26'b01110001010010110000110000 :
  (x[23:13] == 447) ? 26'b01110001010000010011000100 :
  (x[23:13] == 448) ? 26'b01110001001101110101100010 :
  (x[23:13] == 449) ? 26'b01110001001011011000001100 :
  (x[23:13] == 450) ? 26'b01110001001000111010111010 :
  (x[23:13] == 451) ? 26'b01110001000110011101111000 :
  (x[23:13] == 452) ? 26'b01110001000100000000111100 :
  (x[23:13] == 453) ? 26'b01110001000001100100010000 :
  (x[23:13] == 454) ? 26'b01110000111111000111101000 :
  (x[23:13] == 455) ? 26'b01110000111100101011001100 :
  (x[23:13] == 456) ? 26'b01110000111010001110111100 :
  (x[23:13] == 457) ? 26'b01110000110111110010110100 :
  (x[23:13] == 458) ? 26'b01110000110101010110111000 :
  (x[23:13] == 459) ? 26'b01110000110010111011000100 :
  (x[23:13] == 460) ? 26'b01110000110000011111011100 :
  (x[23:13] == 461) ? 26'b01110000101110000011111100 :
  (x[23:13] == 462) ? 26'b01110000101011101000101000 :
  (x[23:13] == 463) ? 26'b01110000101001001101011100 :
  (x[23:13] == 464) ? 26'b01110000100110110010011100 :
  (x[23:13] == 465) ? 26'b01110000100100010111101000 :
  (x[23:13] == 466) ? 26'b01110000100001111100111000 :
  (x[23:13] == 467) ? 26'b01110000011111100010011000 :
  (x[23:13] == 468) ? 26'b01110000011101000111111110 :
  (x[23:13] == 469) ? 26'b01110000011010101101110000 :
  (x[23:13] == 470) ? 26'b01110000011000010011101100 :
  (x[23:13] == 471) ? 26'b01110000010101111001110000 :
  (x[23:13] == 472) ? 26'b01110000010011100000000000 :
  (x[23:13] == 473) ? 26'b01110000010001000110010100 :
  (x[23:13] == 474) ? 26'b01110000001110101100111010 :
  (x[23:13] == 475) ? 26'b01110000001100010011100100 :
  (x[23:13] == 476) ? 26'b01110000001001111010011100 :
  (x[23:13] == 477) ? 26'b01110000000111100001011100 :
  (x[23:13] == 478) ? 26'b01110000000101001000100100 :
  (x[23:13] == 479) ? 26'b01110000000010101111111000 :
  (x[23:13] == 480) ? 26'b01110000000000010111010100 :
  (x[23:13] == 481) ? 26'b01101111111101111110111100 :
  (x[23:13] == 482) ? 26'b01101111111011100110101100 :
  (x[23:13] == 483) ? 26'b01101111111001001110101000 :
  (x[23:13] == 484) ? 26'b01101111110110110110101010 :
  (x[23:13] == 485) ? 26'b01101111110100011110111000 :
  (x[23:13] == 486) ? 26'b01101111110010000111010000 :
  (x[23:13] == 487) ? 26'b01101111101111101111110010 :
  (x[23:13] == 488) ? 26'b01101111101101011000011100 :
  (x[23:13] == 489) ? 26'b01101111101011000001010000 :
  (x[23:13] == 490) ? 26'b01101111101000101010001110 :
  (x[23:13] == 491) ? 26'b01101111100110010011010100 :
  (x[23:13] == 492) ? 26'b01101111100011111100100100 :
  (x[23:13] == 493) ? 26'b01101111100001100110000000 :
  (x[23:13] == 494) ? 26'b01101111011111001111100100 :
  (x[23:13] == 495) ? 26'b01101111011100111001010000 :
  (x[23:13] == 496) ? 26'b01101111011010100011001000 :
  (x[23:13] == 497) ? 26'b01101111011000001101001000 :
  (x[23:13] == 498) ? 26'b01101111010101110111010100 :
  (x[23:13] == 499) ? 26'b01101111010011100001100110 :
  (x[23:13] == 500) ? 26'b01101111010001001100000100 :
  (x[23:13] == 501) ? 26'b01101111001110110110101000 :
  (x[23:13] == 502) ? 26'b01101111001100100001011000 :
  (x[23:13] == 503) ? 26'b01101111001010001100010000 :
  (x[23:13] == 504) ? 26'b01101111000111110111010100 :
  (x[23:13] == 505) ? 26'b01101111000101100010100000 :
  (x[23:13] == 506) ? 26'b01101111000011001101110100 :
  (x[23:13] == 507) ? 26'b01101111000000111001010010 :
  (x[23:13] == 508) ? 26'b01101110111110100100111100 :
  (x[23:13] == 509) ? 26'b01101110111100010000101100 :
  (x[23:13] == 510) ? 26'b01101110111001111100100100 :
  (x[23:13] == 511) ? 26'b01101110110111101000101000 :
  (x[23:13] == 512) ? 26'b01101110110101010100110110 :
  (x[23:13] == 513) ? 26'b01101110110011000001001100 :
  (x[23:13] == 514) ? 26'b01101110110000101101101100 :
  (x[23:13] == 515) ? 26'b01101110101110011010010100 :
  (x[23:13] == 516) ? 26'b01101110101100000111000100 :
  (x[23:13] == 517) ? 26'b01101110101001110100000000 :
  (x[23:13] == 518) ? 26'b01101110100111100001000100 :
  (x[23:13] == 519) ? 26'b01101110100101001110010000 :
  (x[23:13] == 520) ? 26'b01101110100010111011101000 :
  (x[23:13] == 521) ? 26'b01101110100000101001000110 :
  (x[23:13] == 522) ? 26'b01101110011110010110101100 :
  (x[23:13] == 523) ? 26'b01101110011100000100100000 :
  (x[23:13] == 524) ? 26'b01101110011001110010011000 :
  (x[23:13] == 525) ? 26'b01101110010111100000011110 :
  (x[23:13] == 526) ? 26'b01101110010101001110101000 :
  (x[23:13] == 527) ? 26'b01101110010010111101000000 :
  (x[23:13] == 528) ? 26'b01101110010000101011011100 :
  (x[23:13] == 529) ? 26'b01101110001110011010000110 :
  (x[23:13] == 530) ? 26'b01101110001100001000110100 :
  (x[23:13] == 531) ? 26'b01101110001001110111110000 :
  (x[23:13] == 532) ? 26'b01101110000111100110110000 :
  (x[23:13] == 533) ? 26'b01101110000101010101111110 :
  (x[23:13] == 534) ? 26'b01101110000011000101010000 :
  (x[23:13] == 535) ? 26'b01101110000000110100110000 :
  (x[23:13] == 536) ? 26'b01101101111110100100010100 :
  (x[23:13] == 537) ? 26'b01101101111100010100000110 :
  (x[23:13] == 538) ? 26'b01101101111010000011111100 :
  (x[23:13] == 539) ? 26'b01101101110111110011111100 :
  (x[23:13] == 540) ? 26'b01101101110101100100000110 :
  (x[23:13] == 541) ? 26'b01101101110011010100011000 :
  (x[23:13] == 542) ? 26'b01101101110001000100110100 :
  (x[23:13] == 543) ? 26'b01101101101110110101011000 :
  (x[23:13] == 544) ? 26'b01101101101100100110000100 :
  (x[23:13] == 545) ? 26'b01101101101010010110111010 :
  (x[23:13] == 546) ? 26'b01101101101000000111111000 :
  (x[23:13] == 547) ? 26'b01101101100101111001000000 :
  (x[23:13] == 548) ? 26'b01101101100011101010010000 :
  (x[23:13] == 549) ? 26'b01101101100001011011101000 :
  (x[23:13] == 550) ? 26'b01101101011111001101001000 :
  (x[23:13] == 551) ? 26'b01101101011100111110110010 :
  (x[23:13] == 552) ? 26'b01101101011010110000101000 :
  (x[23:13] == 553) ? 26'b01101101011000100010100010 :
  (x[23:13] == 554) ? 26'b01101101010110010100100110 :
  (x[23:13] == 555) ? 26'b01101101010100000110110000 :
  (x[23:13] == 556) ? 26'b01101101010001111001000110 :
  (x[23:13] == 557) ? 26'b01101101001111101011100100 :
  (x[23:13] == 558) ? 26'b01101101001101011110001010 :
  (x[23:13] == 559) ? 26'b01101101001011010000111000 :
  (x[23:13] == 560) ? 26'b01101101001001000011110010 :
  (x[23:13] == 561) ? 26'b01101101000110110110110000 :
  (x[23:13] == 562) ? 26'b01101101000100101001111000 :
  (x[23:13] == 563) ? 26'b01101101000010011101001010 :
  (x[23:13] == 564) ? 26'b01101101000000010000100010 :
  (x[23:13] == 565) ? 26'b01101100111110000100000110 :
  (x[23:13] == 566) ? 26'b01101100111011110111110000 :
  (x[23:13] == 567) ? 26'b01101100111001101011100100 :
  (x[23:13] == 568) ? 26'b01101100110111011111100000 :
  (x[23:13] == 569) ? 26'b01101100110101010011100000 :
  (x[23:13] == 570) ? 26'b01101100110011000111110000 :
  (x[23:13] == 571) ? 26'b01101100110000111100000100 :
  (x[23:13] == 572) ? 26'b01101100101110110000100000 :
  (x[23:13] == 573) ? 26'b01101100101100100101000110 :
  (x[23:13] == 574) ? 26'b01101100101010011001110010 :
  (x[23:13] == 575) ? 26'b01101100101000001110101010 :
  (x[23:13] == 576) ? 26'b01101100100110000011101000 :
  (x[23:13] == 577) ? 26'b01101100100011111000110000 :
  (x[23:13] == 578) ? 26'b01101100100001101110000000 :
  (x[23:13] == 579) ? 26'b01101100011111100011010100 :
  (x[23:13] == 580) ? 26'b01101100011101011000110100 :
  (x[23:13] == 581) ? 26'b01101100011011001110011100 :
  (x[23:13] == 582) ? 26'b01101100011001000100001100 :
  (x[23:13] == 583) ? 26'b01101100010110111010001000 :
  (x[23:13] == 584) ? 26'b01101100010100110000001000 :
  (x[23:13] == 585) ? 26'b01101100010010100110010000 :
  (x[23:13] == 586) ? 26'b01101100010000011100100010 :
  (x[23:13] == 587) ? 26'b01101100001110010010111010 :
  (x[23:13] == 588) ? 26'b01101100001100001001011110 :
  (x[23:13] == 589) ? 26'b01101100001010000000001000 :
  (x[23:13] == 590) ? 26'b01101100000111110110111000 :
  (x[23:13] == 591) ? 26'b01101100000101101101110100 :
  (x[23:13] == 592) ? 26'b01101100000011100100110110 :
  (x[23:13] == 593) ? 26'b01101100000001011100000000 :
  (x[23:13] == 594) ? 26'b01101011111111010011010010 :
  (x[23:13] == 595) ? 26'b01101011111101001010101100 :
  (x[23:13] == 596) ? 26'b01101011111011000010010000 :
  (x[23:13] == 597) ? 26'b01101011111000111001111100 :
  (x[23:13] == 598) ? 26'b01101011110110110001101100 :
  (x[23:13] == 599) ? 26'b01101011110100101001101000 :
  (x[23:13] == 600) ? 26'b01101011110010100001101100 :
  (x[23:13] == 601) ? 26'b01101011110000011001110110 :
  (x[23:13] == 602) ? 26'b01101011101110010010001000 :
  (x[23:13] == 603) ? 26'b01101011101100001010100100 :
  (x[23:13] == 604) ? 26'b01101011101010000011001000 :
  (x[23:13] == 605) ? 26'b01101011100111111011110010 :
  (x[23:13] == 606) ? 26'b01101011100101110100100110 :
  (x[23:13] == 607) ? 26'b01101011100011101101100000 :
  (x[23:13] == 608) ? 26'b01101011100001100110100100 :
  (x[23:13] == 609) ? 26'b01101011011111011111110000 :
  (x[23:13] == 610) ? 26'b01101011011101011001000000 :
  (x[23:13] == 611) ? 26'b01101011011011010010011100 :
  (x[23:13] == 612) ? 26'b01101011011001001100000000 :
  (x[23:13] == 613) ? 26'b01101011010111000101101010 :
  (x[23:13] == 614) ? 26'b01101011010100111111011100 :
  (x[23:13] == 615) ? 26'b01101011010010111001010110 :
  (x[23:13] == 616) ? 26'b01101011010000110011011000 :
  (x[23:13] == 617) ? 26'b01101011001110101101100100 :
  (x[23:13] == 618) ? 26'b01101011001100100111110100 :
  (x[23:13] == 619) ? 26'b01101011001010100010001110 :
  (x[23:13] == 620) ? 26'b01101011001000011100101110 :
  (x[23:13] == 621) ? 26'b01101011000110010111011000 :
  (x[23:13] == 622) ? 26'b01101011000100010010001000 :
  (x[23:13] == 623) ? 26'b01101011000010001101000000 :
  (x[23:13] == 624) ? 26'b01101011000000001000000010 :
  (x[23:13] == 625) ? 26'b01101010111110000011001000 :
  (x[23:13] == 626) ? 26'b01101010111011111110011000 :
  (x[23:13] == 627) ? 26'b01101010111001111001110010 :
  (x[23:13] == 628) ? 26'b01101010110111110101010000 :
  (x[23:13] == 629) ? 26'b01101010110101110000111000 :
  (x[23:13] == 630) ? 26'b01101010110011101100101000 :
  (x[23:13] == 631) ? 26'b01101010110001101000011110 :
  (x[23:13] == 632) ? 26'b01101010101111100100011100 :
  (x[23:13] == 633) ? 26'b01101010101101100000100000 :
  (x[23:13] == 634) ? 26'b01101010101011011100101100 :
  (x[23:13] == 635) ? 26'b01101010101001011001000010 :
  (x[23:13] == 636) ? 26'b01101010100111010101100000 :
  (x[23:13] == 637) ? 26'b01101010100101010010000100 :
  (x[23:13] == 638) ? 26'b01101010100011001110101110 :
  (x[23:13] == 639) ? 26'b01101010100001001011100100 :
  (x[23:13] == 640) ? 26'b01101010011111001000011100 :
  (x[23:13] == 641) ? 26'b01101010011101000101100000 :
  (x[23:13] == 642) ? 26'b01101010011011000010101010 :
  (x[23:13] == 643) ? 26'b01101010011000111111111100 :
  (x[23:13] == 644) ? 26'b01101010010110111101010100 :
  (x[23:13] == 645) ? 26'b01101010010100111010110100 :
  (x[23:13] == 646) ? 26'b01101010010010111000011110 :
  (x[23:13] == 647) ? 26'b01101010010000110110001100 :
  (x[23:13] == 648) ? 26'b01101010001110110100000100 :
  (x[23:13] == 649) ? 26'b01101010001100110010000100 :
  (x[23:13] == 650) ? 26'b01101010001010110000001000 :
  (x[23:13] == 651) ? 26'b01101010001000101110010100 :
  (x[23:13] == 652) ? 26'b01101010000110101100101010 :
  (x[23:13] == 653) ? 26'b01101010000100101011000110 :
  (x[23:13] == 654) ? 26'b01101010000010101001101100 :
  (x[23:13] == 655) ? 26'b01101010000000101000010110 :
  (x[23:13] == 656) ? 26'b01101001111110100111001000 :
  (x[23:13] == 657) ? 26'b01101001111100100110000000 :
  (x[23:13] == 658) ? 26'b01101001111010100101000100 :
  (x[23:13] == 659) ? 26'b01101001111000100100001010 :
  (x[23:13] == 660) ? 26'b01101001110110100011011100 :
  (x[23:13] == 661) ? 26'b01101001110100100010110000 :
  (x[23:13] == 662) ? 26'b01101001110010100010010010 :
  (x[23:13] == 663) ? 26'b01101001110000100001110110 :
  (x[23:13] == 664) ? 26'b01101001101110100001100100 :
  (x[23:13] == 665) ? 26'b01101001101100100001011000 :
  (x[23:13] == 666) ? 26'b01101001101010100001010100 :
  (x[23:13] == 667) ? 26'b01101001101000100001011000 :
  (x[23:13] == 668) ? 26'b01101001100110100001100010 :
  (x[23:13] == 669) ? 26'b01101001100100100001110100 :
  (x[23:13] == 670) ? 26'b01101001100010100010001100 :
  (x[23:13] == 671) ? 26'b01101001100000100010101100 :
  (x[23:13] == 672) ? 26'b01101001011110100011010100 :
  (x[23:13] == 673) ? 26'b01101001011100100100000010 :
  (x[23:13] == 674) ? 26'b01101001011010100100111000 :
  (x[23:13] == 675) ? 26'b01101001011000100101110010 :
  (x[23:13] == 676) ? 26'b01101001010110100110110110 :
  (x[23:13] == 677) ? 26'b01101001010100101000000100 :
  (x[23:13] == 678) ? 26'b01101001010010101001010110 :
  (x[23:13] == 679) ? 26'b01101001010000101010110000 :
  (x[23:13] == 680) ? 26'b01101001001110101100001110 :
  (x[23:13] == 681) ? 26'b01101001001100101101110110 :
  (x[23:13] == 682) ? 26'b01101001001010101111100100 :
  (x[23:13] == 683) ? 26'b01101001001000110001011100 :
  (x[23:13] == 684) ? 26'b01101001000110110011011000 :
  (x[23:13] == 685) ? 26'b01101001000100110101011100 :
  (x[23:13] == 686) ? 26'b01101001000010110111101000 :
  (x[23:13] == 687) ? 26'b01101001000000111001111000 :
  (x[23:13] == 688) ? 26'b01101000111110111100010000 :
  (x[23:13] == 689) ? 26'b01101000111100111110110010 :
  (x[23:13] == 690) ? 26'b01101000111011000001011000 :
  (x[23:13] == 691) ? 26'b01101000111001000100001000 :
  (x[23:13] == 692) ? 26'b01101000110111000111000000 :
  (x[23:13] == 693) ? 26'b01101000110101001001111100 :
  (x[23:13] == 694) ? 26'b01101000110011001100111100 :
  (x[23:13] == 695) ? 26'b01101000110001010000001000 :
  (x[23:13] == 696) ? 26'b01101000101111010011011000 :
  (x[23:13] == 697) ? 26'b01101000101101010110110000 :
  (x[23:13] == 698) ? 26'b01101000101011011010010000 :
  (x[23:13] == 699) ? 26'b01101000101001011101110110 :
  (x[23:13] == 700) ? 26'b01101000100111100001100010 :
  (x[23:13] == 701) ? 26'b01101000100101100101011000 :
  (x[23:13] == 702) ? 26'b01101000100011101001010010 :
  (x[23:13] == 703) ? 26'b01101000100001101101010100 :
  (x[23:13] == 704) ? 26'b01101000011111110001011100 :
  (x[23:13] == 705) ? 26'b01101000011101110101101100 :
  (x[23:13] == 706) ? 26'b01101000011011111010000100 :
  (x[23:13] == 707) ? 26'b01101000011001111110100000 :
  (x[23:13] == 708) ? 26'b01101000011000000011000100 :
  (x[23:13] == 709) ? 26'b01101000010110000111110000 :
  (x[23:13] == 710) ? 26'b01101000010100001100100000 :
  (x[23:13] == 711) ? 26'b01101000010010010001011000 :
  (x[23:13] == 712) ? 26'b01101000010000010110011000 :
  (x[23:13] == 713) ? 26'b01101000001110011011011100 :
  (x[23:13] == 714) ? 26'b01101000001100100000101100 :
  (x[23:13] == 715) ? 26'b01101000001010100101111110 :
  (x[23:13] == 716) ? 26'b01101000001000101011011000 :
  (x[23:13] == 717) ? 26'b01101000000110110000111010 :
  (x[23:13] == 718) ? 26'b01101000000100110110100000 :
  (x[23:13] == 719) ? 26'b01101000000010111100010000 :
  (x[23:13] == 720) ? 26'b01101000000001000010001000 :
  (x[23:13] == 721) ? 26'b01100111111111001000000100 :
  (x[23:13] == 722) ? 26'b01100111111101001110000100 :
  (x[23:13] == 723) ? 26'b01100111111011010100010000 :
  (x[23:13] == 724) ? 26'b01100111111001011010011110 :
  (x[23:13] == 725) ? 26'b01100111110111100000110100 :
  (x[23:13] == 726) ? 26'b01100111110101100111010100 :
  (x[23:13] == 727) ? 26'b01100111110011101101111000 :
  (x[23:13] == 728) ? 26'b01100111110001110100100100 :
  (x[23:13] == 729) ? 26'b01100111101111111011010110 :
  (x[23:13] == 730) ? 26'b01100111101110000010001110 :
  (x[23:13] == 731) ? 26'b01100111101100001001001100 :
  (x[23:13] == 732) ? 26'b01100111101010010000010000 :
  (x[23:13] == 733) ? 26'b01100111101000010111011100 :
  (x[23:13] == 734) ? 26'b01100111100110011110110000 :
  (x[23:13] == 735) ? 26'b01100111100100100110001000 :
  (x[23:13] == 736) ? 26'b01100111100010101101101000 :
  (x[23:13] == 737) ? 26'b01100111100000110101010000 :
  (x[23:13] == 738) ? 26'b01100111011110111100111100 :
  (x[23:13] == 739) ? 26'b01100111011101000100110000 :
  (x[23:13] == 740) ? 26'b01100111011011001100101000 :
  (x[23:13] == 741) ? 26'b01100111011001010100101000 :
  (x[23:13] == 742) ? 26'b01100111010111011100110010 :
  (x[23:13] == 743) ? 26'b01100111010101100100111110 :
  (x[23:13] == 744) ? 26'b01100111010011101101010100 :
  (x[23:13] == 745) ? 26'b01100111010001110101101110 :
  (x[23:13] == 746) ? 26'b01100111001111111110010000 :
  (x[23:13] == 747) ? 26'b01100111001110000110110110 :
  (x[23:13] == 748) ? 26'b01100111001100001111100100 :
  (x[23:13] == 749) ? 26'b01100111001010011000011000 :
  (x[23:13] == 750) ? 26'b01100111001000100001010100 :
  (x[23:13] == 751) ? 26'b01100111000110101010010100 :
  (x[23:13] == 752) ? 26'b01100111000100110011011100 :
  (x[23:13] == 753) ? 26'b01100111000010111100101010 :
  (x[23:13] == 754) ? 26'b01100111000001000110000000 :
  (x[23:13] == 755) ? 26'b01100110111111001111011100 :
  (x[23:13] == 756) ? 26'b01100110111101011000111100 :
  (x[23:13] == 757) ? 26'b01100110111011100010100100 :
  (x[23:13] == 758) ? 26'b01100110111001101100010100 :
  (x[23:13] == 759) ? 26'b01100110110111110110001000 :
  (x[23:13] == 760) ? 26'b01100110110110000000000100 :
  (x[23:13] == 761) ? 26'b01100110110100001010000100 :
  (x[23:13] == 762) ? 26'b01100110110010010100001100 :
  (x[23:13] == 763) ? 26'b01100110110000011110011000 :
  (x[23:13] == 764) ? 26'b01100110101110101000101110 :
  (x[23:13] == 765) ? 26'b01100110101100110011001000 :
  (x[23:13] == 766) ? 26'b01100110101010111101101000 :
  (x[23:13] == 767) ? 26'b01100110101001001000010000 :
  (x[23:13] == 768) ? 26'b01100110100111010010111100 :
  (x[23:13] == 769) ? 26'b01100110100101011101110000 :
  (x[23:13] == 770) ? 26'b01100110100011101000101010 :
  (x[23:13] == 771) ? 26'b01100110100001110011101010 :
  (x[23:13] == 772) ? 26'b01100110011111111110110100 :
  (x[23:13] == 773) ? 26'b01100110011110001010000000 :
  (x[23:13] == 774) ? 26'b01100110011100010101010000 :
  (x[23:13] == 775) ? 26'b01100110011010100000101100 :
  (x[23:13] == 776) ? 26'b01100110011000101100001010 :
  (x[23:13] == 777) ? 26'b01100110010110110111110000 :
  (x[23:13] == 778) ? 26'b01100110010101000011011100 :
  (x[23:13] == 779) ? 26'b01100110010011001111001110 :
  (x[23:13] == 780) ? 26'b01100110010001011011001000 :
  (x[23:13] == 781) ? 26'b01100110001111100111000100 :
  (x[23:13] == 782) ? 26'b01100110001101110011001000 :
  (x[23:13] == 783) ? 26'b01100110001011111111010100 :
  (x[23:13] == 784) ? 26'b01100110001010001011100100 :
  (x[23:13] == 785) ? 26'b01100110001000010111111100 :
  (x[23:13] == 786) ? 26'b01100110000110100100011000 :
  (x[23:13] == 787) ? 26'b01100110000100110000111100 :
  (x[23:13] == 788) ? 26'b01100110000010111101101000 :
  (x[23:13] == 789) ? 26'b01100110000001001010010110 :
  (x[23:13] == 790) ? 26'b01100101111111010111001100 :
  (x[23:13] == 791) ? 26'b01100101111101100100000110 :
  (x[23:13] == 792) ? 26'b01100101111011110001001000 :
  (x[23:13] == 793) ? 26'b01100101111001111110010000 :
  (x[23:13] == 794) ? 26'b01100101111000001011011110 :
  (x[23:13] == 795) ? 26'b01100101110110011000110000 :
  (x[23:13] == 796) ? 26'b01100101110100100110001100 :
  (x[23:13] == 797) ? 26'b01100101110010110011101100 :
  (x[23:13] == 798) ? 26'b01100101110001000001010000 :
  (x[23:13] == 799) ? 26'b01100101101111001111000000 :
  (x[23:13] == 800) ? 26'b01100101101101011100110000 :
  (x[23:13] == 801) ? 26'b01100101101011101010101010 :
  (x[23:13] == 802) ? 26'b01100101101001111000101000 :
  (x[23:13] == 803) ? 26'b01100101101000000110101010 :
  (x[23:13] == 804) ? 26'b01100101100110010100110110 :
  (x[23:13] == 805) ? 26'b01100101100100100011000100 :
  (x[23:13] == 806) ? 26'b01100101100010110001011010 :
  (x[23:13] == 807) ? 26'b01100101100000111111111000 :
  (x[23:13] == 808) ? 26'b01100101011111001110011000 :
  (x[23:13] == 809) ? 26'b01100101011101011101000000 :
  (x[23:13] == 810) ? 26'b01100101011011101011110000 :
  (x[23:13] == 811) ? 26'b01100101011001111010100100 :
  (x[23:13] == 812) ? 26'b01100101011000001001011100 :
  (x[23:13] == 813) ? 26'b01100101010110011000011100 :
  (x[23:13] == 814) ? 26'b01100101010100100111100000 :
  (x[23:13] == 815) ? 26'b01100101010010110110101110 :
  (x[23:13] == 816) ? 26'b01100101010001000110000000 :
  (x[23:13] == 817) ? 26'b01100101001111010101010110 :
  (x[23:13] == 818) ? 26'b01100101001101100100110100 :
  (x[23:13] == 819) ? 26'b01100101001011110100010110 :
  (x[23:13] == 820) ? 26'b01100101001010000100000000 :
  (x[23:13] == 821) ? 26'b01100101001000010011101100 :
  (x[23:13] == 822) ? 26'b01100101000110100011100000 :
  (x[23:13] == 823) ? 26'b01100101000100110011011100 :
  (x[23:13] == 824) ? 26'b01100101000011000011011100 :
  (x[23:13] == 825) ? 26'b01100101000001010011100000 :
  (x[23:13] == 826) ? 26'b01100100111111100011101100 :
  (x[23:13] == 827) ? 26'b01100100111101110011111100 :
  (x[23:13] == 828) ? 26'b01100100111100000100010110 :
  (x[23:13] == 829) ? 26'b01100100111010010100110010 :
  (x[23:13] == 830) ? 26'b01100100111000100101011000 :
  (x[23:13] == 831) ? 26'b01100100110110110110000000 :
  (x[23:13] == 832) ? 26'b01100100110101000110101100 :
  (x[23:13] == 833) ? 26'b01100100110011010111100000 :
  (x[23:13] == 834) ? 26'b01100100110001101000011100 :
  (x[23:13] == 835) ? 26'b01100100101111111001011100 :
  (x[23:13] == 836) ? 26'b01100100101110001010011110 :
  (x[23:13] == 837) ? 26'b01100100101100011011101010 :
  (x[23:13] == 838) ? 26'b01100100101010101100111100 :
  (x[23:13] == 839) ? 26'b01100100101000111110010000 :
  (x[23:13] == 840) ? 26'b01100100100111001111110000 :
  (x[23:13] == 841) ? 26'b01100100100101100001010000 :
  (x[23:13] == 842) ? 26'b01100100100011110010111000 :
  (x[23:13] == 843) ? 26'b01100100100010000100100100 :
  (x[23:13] == 844) ? 26'b01100100100000010110011000 :
  (x[23:13] == 845) ? 26'b01100100011110101000010000 :
  (x[23:13] == 846) ? 26'b01100100011100111010010000 :
  (x[23:13] == 847) ? 26'b01100100011011001100010000 :
  (x[23:13] == 848) ? 26'b01100100011001011110011100 :
  (x[23:13] == 849) ? 26'b01100100010111110000101010 :
  (x[23:13] == 850) ? 26'b01100100010110000010111110 :
  (x[23:13] == 851) ? 26'b01100100010100010101011100 :
  (x[23:13] == 852) ? 26'b01100100010010100111111100 :
  (x[23:13] == 853) ? 26'b01100100010000111010011110 :
  (x[23:13] == 854) ? 26'b01100100001111001101001010 :
  (x[23:13] == 855) ? 26'b01100100001101011111111100 :
  (x[23:13] == 856) ? 26'b01100100001011110010110000 :
  (x[23:13] == 857) ? 26'b01100100001010000101101100 :
  (x[23:13] == 858) ? 26'b01100100001000011000110000 :
  (x[23:13] == 859) ? 26'b01100100000110101011111000 :
  (x[23:13] == 860) ? 26'b01100100000100111111000000 :
  (x[23:13] == 861) ? 26'b01100100000011010010010100 :
  (x[23:13] == 862) ? 26'b01100100000001100101101100 :
  (x[23:13] == 863) ? 26'b01100011111111111001001000 :
  (x[23:13] == 864) ? 26'b01100011111110001100101100 :
  (x[23:13] == 865) ? 26'b01100011111100100000010100 :
  (x[23:13] == 866) ? 26'b01100011111010110100000000 :
  (x[23:13] == 867) ? 26'b01100011111001000111110100 :
  (x[23:13] == 868) ? 26'b01100011110111011011101100 :
  (x[23:13] == 869) ? 26'b01100011110101101111101100 :
  (x[23:13] == 870) ? 26'b01100011110100000011110000 :
  (x[23:13] == 871) ? 26'b01100011110010010111111000 :
  (x[23:13] == 872) ? 26'b01100011110000101100001000 :
  (x[23:13] == 873) ? 26'b01100011101111000000011100 :
  (x[23:13] == 874) ? 26'b01100011101101010100110100 :
  (x[23:13] == 875) ? 26'b01100011101011101001010010 :
  (x[23:13] == 876) ? 26'b01100011101001111101111000 :
  (x[23:13] == 877) ? 26'b01100011101000010010100000 :
  (x[23:13] == 878) ? 26'b01100011100110100111010000 :
  (x[23:13] == 879) ? 26'b01100011100100111100000110 :
  (x[23:13] == 880) ? 26'b01100011100011010001000000 :
  (x[23:13] == 881) ? 26'b01100011100001100101111110 :
  (x[23:13] == 882) ? 26'b01100011011111111011000100 :
  (x[23:13] == 883) ? 26'b01100011011110010000001110 :
  (x[23:13] == 884) ? 26'b01100011011100100101011100 :
  (x[23:13] == 885) ? 26'b01100011011010111010110100 :
  (x[23:13] == 886) ? 26'b01100011011001010000001100 :
  (x[23:13] == 887) ? 26'b01100011010111100101101010 :
  (x[23:13] == 888) ? 26'b01100011010101111011010000 :
  (x[23:13] == 889) ? 26'b01100011010100010000111100 :
  (x[23:13] == 890) ? 26'b01100011010010100110101100 :
  (x[23:13] == 891) ? 26'b01100011010000111100100000 :
  (x[23:13] == 892) ? 26'b01100011001111010010011100 :
  (x[23:13] == 893) ? 26'b01100011001101101000011000 :
  (x[23:13] == 894) ? 26'b01100011001011111110011100 :
  (x[23:13] == 895) ? 26'b01100011001010010100101000 :
  (x[23:13] == 896) ? 26'b01100011001000101010111000 :
  (x[23:13] == 897) ? 26'b01100011000111000001001100 :
  (x[23:13] == 898) ? 26'b01100011000101010111100110 :
  (x[23:13] == 899) ? 26'b01100011000011101110000100 :
  (x[23:13] == 900) ? 26'b01100011000010000100101010 :
  (x[23:13] == 901) ? 26'b01100011000000011011010100 :
  (x[23:13] == 902) ? 26'b01100010111110110010000100 :
  (x[23:13] == 903) ? 26'b01100010111101001000111000 :
  (x[23:13] == 904) ? 26'b01100010111011011111110000 :
  (x[23:13] == 905) ? 26'b01100010111001110110110000 :
  (x[23:13] == 906) ? 26'b01100010111000001101110100 :
  (x[23:13] == 907) ? 26'b01100010110110100100111100 :
  (x[23:13] == 908) ? 26'b01100010110100111100001100 :
  (x[23:13] == 909) ? 26'b01100010110011010011011110 :
  (x[23:13] == 910) ? 26'b01100010110001101010111000 :
  (x[23:13] == 911) ? 26'b01100010110000000010011000 :
  (x[23:13] == 912) ? 26'b01100010101110011001111000 :
  (x[23:13] == 913) ? 26'b01100010101100110001100010 :
  (x[23:13] == 914) ? 26'b01100010101011001001010000 :
  (x[23:13] == 915) ? 26'b01100010101001100001000010 :
  (x[23:13] == 916) ? 26'b01100010100111111000111100 :
  (x[23:13] == 917) ? 26'b01100010100110010000111000 :
  (x[23:13] == 918) ? 26'b01100010100100101000111000 :
  (x[23:13] == 919) ? 26'b01100010100011000001000000 :
  (x[23:13] == 920) ? 26'b01100010100001011001001100 :
  (x[23:13] == 921) ? 26'b01100010011111110001011100 :
  (x[23:13] == 922) ? 26'b01100010011110001001110100 :
  (x[23:13] == 923) ? 26'b01100010011100100010010000 :
  (x[23:13] == 924) ? 26'b01100010011010111010110000 :
  (x[23:13] == 925) ? 26'b01100010011001010011011000 :
  (x[23:13] == 926) ? 26'b01100010010111101100000100 :
  (x[23:13] == 927) ? 26'b01100010010110000100110010 :
  (x[23:13] == 928) ? 26'b01100010010100011101101000 :
  (x[23:13] == 929) ? 26'b01100010010010110110100010 :
  (x[23:13] == 930) ? 26'b01100010010001001111100100 :
  (x[23:13] == 931) ? 26'b01100010001111101000101000 :
  (x[23:13] == 932) ? 26'b01100010001110000001101110 :
  (x[23:13] == 933) ? 26'b01100010001100011010111110 :
  (x[23:13] == 934) ? 26'b01100010001010110100010000 :
  (x[23:13] == 935) ? 26'b01100010001001001101101010 :
  (x[23:13] == 936) ? 26'b01100010000111100111001000 :
  (x[23:13] == 937) ? 26'b01100010000110000000101100 :
  (x[23:13] == 938) ? 26'b01100010000100011010010100 :
  (x[23:13] == 939) ? 26'b01100010000010110011111110 :
  (x[23:13] == 940) ? 26'b01100010000001001101110000 :
  (x[23:13] == 941) ? 26'b01100001111111100111100110 :
  (x[23:13] == 942) ? 26'b01100001111110000001100100 :
  (x[23:13] == 943) ? 26'b01100001111100011011100100 :
  (x[23:13] == 944) ? 26'b01100001111010110101101000 :
  (x[23:13] == 945) ? 26'b01100001111001001111110010 :
  (x[23:13] == 946) ? 26'b01100001110111101010000100 :
  (x[23:13] == 947) ? 26'b01100001110110000100010110 :
  (x[23:13] == 948) ? 26'b01100001110100011110110000 :
  (x[23:13] == 949) ? 26'b01100001110010111001010000 :
  (x[23:13] == 950) ? 26'b01100001110001010011110100 :
  (x[23:13] == 951) ? 26'b01100001101111101110011010 :
  (x[23:13] == 952) ? 26'b01100001101110001001001000 :
  (x[23:13] == 953) ? 26'b01100001101100100011111010 :
  (x[23:13] == 954) ? 26'b01100001101010111110110000 :
  (x[23:13] == 955) ? 26'b01100001101001011001101100 :
  (x[23:13] == 956) ? 26'b01100001100111110100101110 :
  (x[23:13] == 957) ? 26'b01100001100110001111110100 :
  (x[23:13] == 958) ? 26'b01100001100100101010111110 :
  (x[23:13] == 959) ? 26'b01100001100011000110001100 :
  (x[23:13] == 960) ? 26'b01100001100001100001100100 :
  (x[23:13] == 961) ? 26'b01100001011111111100111010 :
  (x[23:13] == 962) ? 26'b01100001011110011000011010 :
  (x[23:13] == 963) ? 26'b01100001011100110011111100 :
  (x[23:13] == 964) ? 26'b01100001011011001111100100 :
  (x[23:13] == 965) ? 26'b01100001011001101011010000 :
  (x[23:13] == 966) ? 26'b01100001011000000111000000 :
  (x[23:13] == 967) ? 26'b01100001010110100010111000 :
  (x[23:13] == 968) ? 26'b01100001010100111110110100 :
  (x[23:13] == 969) ? 26'b01100001010011011010110010 :
  (x[23:13] == 970) ? 26'b01100001010001110110111000 :
  (x[23:13] == 971) ? 26'b01100001010000010011000000 :
  (x[23:13] == 972) ? 26'b01100001001110101111010000 :
  (x[23:13] == 973) ? 26'b01100001001101001011100100 :
  (x[23:13] == 974) ? 26'b01100001001011100111111100 :
  (x[23:13] == 975) ? 26'b01100001001010000100011000 :
  (x[23:13] == 976) ? 26'b01100001001000100000111010 :
  (x[23:13] == 977) ? 26'b01100001000110111101100000 :
  (x[23:13] == 978) ? 26'b01100001000101011010001010 :
  (x[23:13] == 979) ? 26'b01100001000011110110111100 :
  (x[23:13] == 980) ? 26'b01100001000010010011110000 :
  (x[23:13] == 981) ? 26'b01100001000000110000101000 :
  (x[23:13] == 982) ? 26'b01100000111111001101100110 :
  (x[23:13] == 983) ? 26'b01100000111101101010101000 :
  (x[23:13] == 984) ? 26'b01100000111100000111110000 :
  (x[23:13] == 985) ? 26'b01100000111010100100111100 :
  (x[23:13] == 986) ? 26'b01100000111001000010001100 :
  (x[23:13] == 987) ? 26'b01100000110111011111100010 :
  (x[23:13] == 988) ? 26'b01100000110101111100111100 :
  (x[23:13] == 989) ? 26'b01100000110100011010011100 :
  (x[23:13] == 990) ? 26'b01100000110010111000000000 :
  (x[23:13] == 991) ? 26'b01100000110001010101101000 :
  (x[23:13] == 992) ? 26'b01100000101111110011010110 :
  (x[23:13] == 993) ? 26'b01100000101110010001000110 :
  (x[23:13] == 994) ? 26'b01100000101100101111000000 :
  (x[23:13] == 995) ? 26'b01100000101011001100111000 :
  (x[23:13] == 996) ? 26'b01100000101001101010111010 :
  (x[23:13] == 997) ? 26'b01100000101000001000111100 :
  (x[23:13] == 998) ? 26'b01100000100110100111001000 :
  (x[23:13] == 999) ? 26'b01100000100101000101010100 :
  (x[23:13] == 1000) ? 26'b01100000100011100011100110 :
  (x[23:13] == 1001) ? 26'b01100000100010000001111100 :
  (x[23:13] == 1002) ? 26'b01100000100000100000011010 :
  (x[23:13] == 1003) ? 26'b01100000011110111110111010 :
  (x[23:13] == 1004) ? 26'b01100000011101011101011100 :
  (x[23:13] == 1005) ? 26'b01100000011011111100001000 :
  (x[23:13] == 1006) ? 26'b01100000011010011010110100 :
  (x[23:13] == 1007) ? 26'b01100000011000111001101010 :
  (x[23:13] == 1008) ? 26'b01100000010111011000100000 :
  (x[23:13] == 1009) ? 26'b01100000010101110111011100 :
  (x[23:13] == 1010) ? 26'b01100000010100010110011100 :
  (x[23:13] == 1011) ? 26'b01100000010010110101100010 :
  (x[23:13] == 1012) ? 26'b01100000010001010100101100 :
  (x[23:13] == 1013) ? 26'b01100000001111110011111000 :
  (x[23:13] == 1014) ? 26'b01100000001110010011001100 :
  (x[23:13] == 1015) ? 26'b01100000001100110010100010 :
  (x[23:13] == 1016) ? 26'b01100000001011010001111110 :
  (x[23:13] == 1017) ? 26'b01100000001001110001100000 :
  (x[23:13] == 1018) ? 26'b01100000001000010001000100 :
  (x[23:13] == 1019) ? 26'b01100000000110110000101100 :
  (x[23:13] == 1020) ? 26'b01100000000101010000011100 :
  (x[23:13] == 1021) ? 26'b01100000000011110000010000 :
  (x[23:13] == 1022) ? 26'b01100000000010010000000110 :
  (x[23:13] == 1023) ? 26'b01100000000000110000000000 :
  (x[23:13] == 1024) ? 26'b10111111111101000000000100 :
  (x[23:13] == 1025) ? 26'b10111111110111000000101000 :
  (x[23:13] == 1026) ? 26'b10111111110001000001110000 :
  (x[23:13] == 1027) ? 26'b10111111101011000011011100 :
  (x[23:13] == 1028) ? 26'b10111111100101000101101100 :
  (x[23:13] == 1029) ? 26'b10111111011111001000100000 :
  (x[23:13] == 1030) ? 26'b10111111011001001011110100 :
  (x[23:13] == 1031) ? 26'b10111111010011001111101100 :
  (x[23:13] == 1032) ? 26'b10111111001101010100001100 :
  (x[23:13] == 1033) ? 26'b10111111000111011001001100 :
  (x[23:13] == 1034) ? 26'b10111111000001011110110000 :
  (x[23:13] == 1035) ? 26'b10111110111011100100111000 :
  (x[23:13] == 1036) ? 26'b10111110110101101011100000 :
  (x[23:13] == 1037) ? 26'b10111110101111110010110000 :
  (x[23:13] == 1038) ? 26'b10111110101001111010011100 :
  (x[23:13] == 1039) ? 26'b10111110100100000010110000 :
  (x[23:13] == 1040) ? 26'b10111110011110001011100100 :
  (x[23:13] == 1041) ? 26'b10111110011000010100111100 :
  (x[23:13] == 1042) ? 26'b10111110010010011110110100 :
  (x[23:13] == 1043) ? 26'b10111110001100101001010000 :
  (x[23:13] == 1044) ? 26'b10111110000110110100010000 :
  (x[23:13] == 1045) ? 26'b10111110000000111111110000 :
  (x[23:13] == 1046) ? 26'b10111101111011001011110100 :
  (x[23:13] == 1047) ? 26'b10111101110101011000011000 :
  (x[23:13] == 1048) ? 26'b10111101101111100101100000 :
  (x[23:13] == 1049) ? 26'b10111101101001110011001000 :
  (x[23:13] == 1050) ? 26'b10111101100100000001011000 :
  (x[23:13] == 1051) ? 26'b10111101011110010000000000 :
  (x[23:13] == 1052) ? 26'b10111101011000011111010000 :
  (x[23:13] == 1053) ? 26'b10111101010010101111000000 :
  (x[23:13] == 1054) ? 26'b10111101001100111111010000 :
  (x[23:13] == 1055) ? 26'b10111101000111010000001000 :
  (x[23:13] == 1056) ? 26'b10111101000001100001011000 :
  (x[23:13] == 1057) ? 26'b10111100111011110011010000 :
  (x[23:13] == 1058) ? 26'b10111100110110000101101000 :
  (x[23:13] == 1059) ? 26'b10111100110000011000100000 :
  (x[23:13] == 1060) ? 26'b10111100101010101011111000 :
  (x[23:13] == 1061) ? 26'b10111100100100111111110100 :
  (x[23:13] == 1062) ? 26'b10111100011111010100010000 :
  (x[23:13] == 1063) ? 26'b10111100011001101001001000 :
  (x[23:13] == 1064) ? 26'b10111100010011111110101000 :
  (x[23:13] == 1065) ? 26'b10111100001110010100100100 :
  (x[23:13] == 1066) ? 26'b10111100001000101011000100 :
  (x[23:13] == 1067) ? 26'b10111100000011000010000000 :
  (x[23:13] == 1068) ? 26'b10111011111101011001100000 :
  (x[23:13] == 1069) ? 26'b10111011110111110001100000 :
  (x[23:13] == 1070) ? 26'b10111011110010001010000000 :
  (x[23:13] == 1071) ? 26'b10111011101100100011000000 :
  (x[23:13] == 1072) ? 26'b10111011100110111100100000 :
  (x[23:13] == 1073) ? 26'b10111011100001010110100000 :
  (x[23:13] == 1074) ? 26'b10111011011011110001000000 :
  (x[23:13] == 1075) ? 26'b10111011010110001100000000 :
  (x[23:13] == 1076) ? 26'b10111011010000100111100000 :
  (x[23:13] == 1077) ? 26'b10111011001011000011100000 :
  (x[23:13] == 1078) ? 26'b10111011000101100000000000 :
  (x[23:13] == 1079) ? 26'b10111010111111111101000000 :
  (x[23:13] == 1080) ? 26'b10111010111010011010011100 :
  (x[23:13] == 1081) ? 26'b10111010110100111000011100 :
  (x[23:13] == 1082) ? 26'b10111010101111010110111000 :
  (x[23:13] == 1083) ? 26'b10111010101001110101110100 :
  (x[23:13] == 1084) ? 26'b10111010100100010101010000 :
  (x[23:13] == 1085) ? 26'b10111010011110110101001000 :
  (x[23:13] == 1086) ? 26'b10111010011001010101101000 :
  (x[23:13] == 1087) ? 26'b10111010010011110110100000 :
  (x[23:13] == 1088) ? 26'b10111010001110010111111000 :
  (x[23:13] == 1089) ? 26'b10111010001000111001110000 :
  (x[23:13] == 1090) ? 26'b10111010000011011100000100 :
  (x[23:13] == 1091) ? 26'b10111001111101111110111000 :
  (x[23:13] == 1092) ? 26'b10111001111000100010001100 :
  (x[23:13] == 1093) ? 26'b10111001110011000110000000 :
  (x[23:13] == 1094) ? 26'b10111001101101101010010000 :
  (x[23:13] == 1095) ? 26'b10111001101000001110111100 :
  (x[23:13] == 1096) ? 26'b10111001100010110100001100 :
  (x[23:13] == 1097) ? 26'b10111001011101011001111000 :
  (x[23:13] == 1098) ? 26'b10111001011000000000000000 :
  (x[23:13] == 1099) ? 26'b10111001010010100110101000 :
  (x[23:13] == 1100) ? 26'b10111001001101001101110000 :
  (x[23:13] == 1101) ? 26'b10111001000111110101011000 :
  (x[23:13] == 1102) ? 26'b10111001000010011101011000 :
  (x[23:13] == 1103) ? 26'b10111000111101000101111000 :
  (x[23:13] == 1104) ? 26'b10111000110111101110111000 :
  (x[23:13] == 1105) ? 26'b10111000110010011000010000 :
  (x[23:13] == 1106) ? 26'b10111000101101000010001100 :
  (x[23:13] == 1107) ? 26'b10111000100111101100100100 :
  (x[23:13] == 1108) ? 26'b10111000100010010111011000 :
  (x[23:13] == 1109) ? 26'b10111000011101000010101100 :
  (x[23:13] == 1110) ? 26'b10111000010111101110011000 :
  (x[23:13] == 1111) ? 26'b10111000010010011010101000 :
  (x[23:13] == 1112) ? 26'b10111000001101000111010000 :
  (x[23:13] == 1113) ? 26'b10111000000111110100011100 :
  (x[23:13] == 1114) ? 26'b10111000000010100010000000 :
  (x[23:13] == 1115) ? 26'b10110111111101010000000100 :
  (x[23:13] == 1116) ? 26'b10110111110111111110100100 :
  (x[23:13] == 1117) ? 26'b10110111110010101101100000 :
  (x[23:13] == 1118) ? 26'b10110111101101011100111000 :
  (x[23:13] == 1119) ? 26'b10110111101000001100110000 :
  (x[23:13] == 1120) ? 26'b10110111100010111101000000 :
  (x[23:13] == 1121) ? 26'b10110111011101101101110000 :
  (x[23:13] == 1122) ? 26'b10110111011000011111000000 :
  (x[23:13] == 1123) ? 26'b10110111010011010000101000 :
  (x[23:13] == 1124) ? 26'b10110111001110000010101100 :
  (x[23:13] == 1125) ? 26'b10110111001000110101010000 :
  (x[23:13] == 1126) ? 26'b10110111000011101000010000 :
  (x[23:13] == 1127) ? 26'b10110110111110011011101000 :
  (x[23:13] == 1128) ? 26'b10110110111001001111100000 :
  (x[23:13] == 1129) ? 26'b10110110110100000011110100 :
  (x[23:13] == 1130) ? 26'b10110110101110111000100000 :
  (x[23:13] == 1131) ? 26'b10110110101001101101110000 :
  (x[23:13] == 1132) ? 26'b10110110100100100011011000 :
  (x[23:13] == 1133) ? 26'b10110110011111011001011000 :
  (x[23:13] == 1134) ? 26'b10110110011010001111111100 :
  (x[23:13] == 1135) ? 26'b10110110010101000110110100 :
  (x[23:13] == 1136) ? 26'b10110110001111111110001100 :
  (x[23:13] == 1137) ? 26'b10110110001010110110000000 :
  (x[23:13] == 1138) ? 26'b10110110000101101110001100 :
  (x[23:13] == 1139) ? 26'b10110110000000100110111000 :
  (x[23:13] == 1140) ? 26'b10110101111011100000000000 :
  (x[23:13] == 1141) ? 26'b10110101110110011001100000 :
  (x[23:13] == 1142) ? 26'b10110101110001010011100000 :
  (x[23:13] == 1143) ? 26'b10110101101100001101110100 :
  (x[23:13] == 1144) ? 26'b10110101100111001000101000 :
  (x[23:13] == 1145) ? 26'b10110101100010000011111000 :
  (x[23:13] == 1146) ? 26'b10110101011100111111100000 :
  (x[23:13] == 1147) ? 26'b10110101010111111011101000 :
  (x[23:13] == 1148) ? 26'b10110101010010111000001000 :
  (x[23:13] == 1149) ? 26'b10110101001101110101000000 :
  (x[23:13] == 1150) ? 26'b10110101001000110010011000 :
  (x[23:13] == 1151) ? 26'b10110101000011110000001100 :
  (x[23:13] == 1152) ? 26'b10110100111110101110010100 :
  (x[23:13] == 1153) ? 26'b10110100111001101100111100 :
  (x[23:13] == 1154) ? 26'b10110100110100101100000000 :
  (x[23:13] == 1155) ? 26'b10110100101111101011011100 :
  (x[23:13] == 1156) ? 26'b10110100101010101011010000 :
  (x[23:13] == 1157) ? 26'b10110100100101101011100000 :
  (x[23:13] == 1158) ? 26'b10110100100000101100010000 :
  (x[23:13] == 1159) ? 26'b10110100011011101101010100 :
  (x[23:13] == 1160) ? 26'b10110100010110101110111000 :
  (x[23:13] == 1161) ? 26'b10110100010001110000110000 :
  (x[23:13] == 1162) ? 26'b10110100001100110011001000 :
  (x[23:13] == 1163) ? 26'b10110100000111110101111000 :
  (x[23:13] == 1164) ? 26'b10110100000010111001000000 :
  (x[23:13] == 1165) ? 26'b10110011111101111100100100 :
  (x[23:13] == 1166) ? 26'b10110011111001000000100000 :
  (x[23:13] == 1167) ? 26'b10110011110100000100111000 :
  (x[23:13] == 1168) ? 26'b10110011101111001001101100 :
  (x[23:13] == 1169) ? 26'b10110011101010001110110100 :
  (x[23:13] == 1170) ? 26'b10110011100101010100011100 :
  (x[23:13] == 1171) ? 26'b10110011100000011010011100 :
  (x[23:13] == 1172) ? 26'b10110011011011100000110100 :
  (x[23:13] == 1173) ? 26'b10110011010110100111101000 :
  (x[23:13] == 1174) ? 26'b10110011010001101110110100 :
  (x[23:13] == 1175) ? 26'b10110011001100110110011000 :
  (x[23:13] == 1176) ? 26'b10110011000111111110011000 :
  (x[23:13] == 1177) ? 26'b10110011000011000110110000 :
  (x[23:13] == 1178) ? 26'b10110010111110001111100100 :
  (x[23:13] == 1179) ? 26'b10110010111001011000110000 :
  (x[23:13] == 1180) ? 26'b10110010110100100010010000 :
  (x[23:13] == 1181) ? 26'b10110010101111101100010000 :
  (x[23:13] == 1182) ? 26'b10110010101010110110101000 :
  (x[23:13] == 1183) ? 26'b10110010100110000001011000 :
  (x[23:13] == 1184) ? 26'b10110010100001001100100100 :
  (x[23:13] == 1185) ? 26'b10110010011100011000000100 :
  (x[23:13] == 1186) ? 26'b10110010010111100100000000 :
  (x[23:13] == 1187) ? 26'b10110010010010110000010100 :
  (x[23:13] == 1188) ? 26'b10110010001101111101000000 :
  (x[23:13] == 1189) ? 26'b10110010001001001010001000 :
  (x[23:13] == 1190) ? 26'b10110010000100010111101000 :
  (x[23:13] == 1191) ? 26'b10110001111111100101011100 :
  (x[23:13] == 1192) ? 26'b10110001111010110011101100 :
  (x[23:13] == 1193) ? 26'b10110001110110000010011000 :
  (x[23:13] == 1194) ? 26'b10110001110001010001010100 :
  (x[23:13] == 1195) ? 26'b10110001101100100000110000 :
  (x[23:13] == 1196) ? 26'b10110001100111110000100000 :
  (x[23:13] == 1197) ? 26'b10110001100011000000101100 :
  (x[23:13] == 1198) ? 26'b10110001011110010001010000 :
  (x[23:13] == 1199) ? 26'b10110001011001100010001000 :
  (x[23:13] == 1200) ? 26'b10110001010100110011100000 :
  (x[23:13] == 1201) ? 26'b10110001010000000101001000 :
  (x[23:13] == 1202) ? 26'b10110001001011010111010000 :
  (x[23:13] == 1203) ? 26'b10110001000110101001101000 :
  (x[23:13] == 1204) ? 26'b10110001000001111100011100 :
  (x[23:13] == 1205) ? 26'b10110000111101001111101000 :
  (x[23:13] == 1206) ? 26'b10110000111000100011001100 :
  (x[23:13] == 1207) ? 26'b10110000110011110111001000 :
  (x[23:13] == 1208) ? 26'b10110000101111001011011100 :
  (x[23:13] == 1209) ? 26'b10110000101010100000000100 :
  (x[23:13] == 1210) ? 26'b10110000100101110101001000 :
  (x[23:13] == 1211) ? 26'b10110000100001001010100100 :
  (x[23:13] == 1212) ? 26'b10110000011100100000011000 :
  (x[23:13] == 1213) ? 26'b10110000010111110110100000 :
  (x[23:13] == 1214) ? 26'b10110000010011001101000000 :
  (x[23:13] == 1215) ? 26'b10110000001110100011111100 :
  (x[23:13] == 1216) ? 26'b10110000001001111011001100 :
  (x[23:13] == 1217) ? 26'b10110000000101010010110000 :
  (x[23:13] == 1218) ? 26'b10110000000000101010110000 :
  (x[23:13] == 1219) ? 26'b10101111111100000011001000 :
  (x[23:13] == 1220) ? 26'b10101111110111011011111000 :
  (x[23:13] == 1221) ? 26'b10101111110010110100111100 :
  (x[23:13] == 1222) ? 26'b10101111101110001110011000 :
  (x[23:13] == 1223) ? 26'b10101111101001101000001100 :
  (x[23:13] == 1224) ? 26'b10101111100101000010010100 :
  (x[23:13] == 1225) ? 26'b10101111100000011100110100 :
  (x[23:13] == 1226) ? 26'b10101111011011110111110000 :
  (x[23:13] == 1227) ? 26'b10101111010111010011000000 :
  (x[23:13] == 1228) ? 26'b10101111010010101110100100 :
  (x[23:13] == 1229) ? 26'b10101111001110001010100000 :
  (x[23:13] == 1230) ? 26'b10101111001001100110111000 :
  (x[23:13] == 1231) ? 26'b10101111000101000011100000 :
  (x[23:13] == 1232) ? 26'b10101111000000100000100000 :
  (x[23:13] == 1233) ? 26'b10101110111011111101111000 :
  (x[23:13] == 1234) ? 26'b10101110110111011011101000 :
  (x[23:13] == 1235) ? 26'b10101110110010111001101100 :
  (x[23:13] == 1236) ? 26'b10101110101110011000001000 :
  (x[23:13] == 1237) ? 26'b10101110101001110110111000 :
  (x[23:13] == 1238) ? 26'b10101110100101010110000000 :
  (x[23:13] == 1239) ? 26'b10101110100000110101100000 :
  (x[23:13] == 1240) ? 26'b10101110011100010101011000 :
  (x[23:13] == 1241) ? 26'b10101110010111110101100000 :
  (x[23:13] == 1242) ? 26'b10101110010011010110000100 :
  (x[23:13] == 1243) ? 26'b10101110001110110110111000 :
  (x[23:13] == 1244) ? 26'b10101110001010011000001000 :
  (x[23:13] == 1245) ? 26'b10101110000101111001110000 :
  (x[23:13] == 1246) ? 26'b10101110000001011011101000 :
  (x[23:13] == 1247) ? 26'b10101101111100111101111000 :
  (x[23:13] == 1248) ? 26'b10101101111000100000100000 :
  (x[23:13] == 1249) ? 26'b10101101110100000011011000 :
  (x[23:13] == 1250) ? 26'b10101101101111100110101000 :
  (x[23:13] == 1251) ? 26'b10101101101011001010010100 :
  (x[23:13] == 1252) ? 26'b10101101100110101110010000 :
  (x[23:13] == 1253) ? 26'b10101101100010010010100100 :
  (x[23:13] == 1254) ? 26'b10101101011101110111001100 :
  (x[23:13] == 1255) ? 26'b10101101011001011100001100 :
  (x[23:13] == 1256) ? 26'b10101101010101000001100000 :
  (x[23:13] == 1257) ? 26'b10101101010000100111001000 :
  (x[23:13] == 1258) ? 26'b10101101001100001101001000 :
  (x[23:13] == 1259) ? 26'b10101101000111110011100000 :
  (x[23:13] == 1260) ? 26'b10101101000011011010001000 :
  (x[23:13] == 1261) ? 26'b10101100111111000001001000 :
  (x[23:13] == 1262) ? 26'b10101100111010101000100000 :
  (x[23:13] == 1263) ? 26'b10101100110110010000001000 :
  (x[23:13] == 1264) ? 26'b10101100110001111000001000 :
  (x[23:13] == 1265) ? 26'b10101100101101100000100000 :
  (x[23:13] == 1266) ? 26'b10101100101001001001001000 :
  (x[23:13] == 1267) ? 26'b10101100100100110010001000 :
  (x[23:13] == 1268) ? 26'b10101100100000011011100000 :
  (x[23:13] == 1269) ? 26'b10101100011100000101000100 :
  (x[23:13] == 1270) ? 26'b10101100010111101111000100 :
  (x[23:13] == 1271) ? 26'b10101100010011011001011000 :
  (x[23:13] == 1272) ? 26'b10101100001111000100000000 :
  (x[23:13] == 1273) ? 26'b10101100001010101111000000 :
  (x[23:13] == 1274) ? 26'b10101100000110011010010000 :
  (x[23:13] == 1275) ? 26'b10101100000010000101111000 :
  (x[23:13] == 1276) ? 26'b10101011111101110001110100 :
  (x[23:13] == 1277) ? 26'b10101011111001011110001000 :
  (x[23:13] == 1278) ? 26'b10101011110101001010101000 :
  (x[23:13] == 1279) ? 26'b10101011110000110111101000 :
  (x[23:13] == 1280) ? 26'b10101011101100100100110100 :
  (x[23:13] == 1281) ? 26'b10101011101000010010011000 :
  (x[23:13] == 1282) ? 26'b10101011100100000000010000 :
  (x[23:13] == 1283) ? 26'b10101011011111101110011100 :
  (x[23:13] == 1284) ? 26'b10101011011011011101000000 :
  (x[23:13] == 1285) ? 26'b10101011010111001011110000 :
  (x[23:13] == 1286) ? 26'b10101011010010111011000000 :
  (x[23:13] == 1287) ? 26'b10101011001110101010011100 :
  (x[23:13] == 1288) ? 26'b10101011001010011010001100 :
  (x[23:13] == 1289) ? 26'b10101011000110001010010100 :
  (x[23:13] == 1290) ? 26'b10101011000001111010110000 :
  (x[23:13] == 1291) ? 26'b10101010111101101011011100 :
  (x[23:13] == 1292) ? 26'b10101010111001011100100000 :
  (x[23:13] == 1293) ? 26'b10101010110101001101111000 :
  (x[23:13] == 1294) ? 26'b10101010110000111111100100 :
  (x[23:13] == 1295) ? 26'b10101010101100110001100000 :
  (x[23:13] == 1296) ? 26'b10101010101000100011111000 :
  (x[23:13] == 1297) ? 26'b10101010100100010110100000 :
  (x[23:13] == 1298) ? 26'b10101010100000001001011000 :
  (x[23:13] == 1299) ? 26'b10101010011011111100101000 :
  (x[23:13] == 1300) ? 26'b10101010010111110000001100 :
  (x[23:13] == 1301) ? 26'b10101010010011100100000100 :
  (x[23:13] == 1302) ? 26'b10101010001111011000001100 :
  (x[23:13] == 1303) ? 26'b10101010001011001100101100 :
  (x[23:13] == 1304) ? 26'b10101010000111000001011100 :
  (x[23:13] == 1305) ? 26'b10101010000010110110100100 :
  (x[23:13] == 1306) ? 26'b10101001111110101100000000 :
  (x[23:13] == 1307) ? 26'b10101001111010100001101100 :
  (x[23:13] == 1308) ? 26'b10101001110110010111101000 :
  (x[23:13] == 1309) ? 26'b10101001110010001110000000 :
  (x[23:13] == 1310) ? 26'b10101001101110000100101000 :
  (x[23:13] == 1311) ? 26'b10101001101001111011100000 :
  (x[23:13] == 1312) ? 26'b10101001100101110010110000 :
  (x[23:13] == 1313) ? 26'b10101001100001101010010000 :
  (x[23:13] == 1314) ? 26'b10101001011101100010000100 :
  (x[23:13] == 1315) ? 26'b10101001011001011010010000 :
  (x[23:13] == 1316) ? 26'b10101001010101010010101000 :
  (x[23:13] == 1317) ? 26'b10101001010001001011011000 :
  (x[23:13] == 1318) ? 26'b10101001001101000100011100 :
  (x[23:13] == 1319) ? 26'b10101001001000111101110000 :
  (x[23:13] == 1320) ? 26'b10101001000100110111011000 :
  (x[23:13] == 1321) ? 26'b10101001000000110001010100 :
  (x[23:13] == 1322) ? 26'b10101000111100101011100000 :
  (x[23:13] == 1323) ? 26'b10101000111000100110000000 :
  (x[23:13] == 1324) ? 26'b10101000110100100000111000 :
  (x[23:13] == 1325) ? 26'b10101000110000011011111100 :
  (x[23:13] == 1326) ? 26'b10101000101100010111011000 :
  (x[23:13] == 1327) ? 26'b10101000101000010011000100 :
  (x[23:13] == 1328) ? 26'b10101000100100001111000100 :
  (x[23:13] == 1329) ? 26'b10101000100000001011010100 :
  (x[23:13] == 1330) ? 26'b10101000011100000111111000 :
  (x[23:13] == 1331) ? 26'b10101000011000000100110000 :
  (x[23:13] == 1332) ? 26'b10101000010100000001111100 :
  (x[23:13] == 1333) ? 26'b10101000001111111111011100 :
  (x[23:13] == 1334) ? 26'b10101000001011111101001000 :
  (x[23:13] == 1335) ? 26'b10101000000111111011001100 :
  (x[23:13] == 1336) ? 26'b10101000000011111001100000 :
  (x[23:13] == 1337) ? 26'b10100111111111111000001000 :
  (x[23:13] == 1338) ? 26'b10100111111011110111000000 :
  (x[23:13] == 1339) ? 26'b10100111110111110110010000 :
  (x[23:13] == 1340) ? 26'b10100111110011110101101100 :
  (x[23:13] == 1341) ? 26'b10100111101111110101100000 :
  (x[23:13] == 1342) ? 26'b10100111101011110101100000 :
  (x[23:13] == 1343) ? 26'b10100111100111110101111000 :
  (x[23:13] == 1344) ? 26'b10100111100011110110011100 :
  (x[23:13] == 1345) ? 26'b10100111011111110111011000 :
  (x[23:13] == 1346) ? 26'b10100111011011111000101000 :
  (x[23:13] == 1347) ? 26'b10100111010111111010000100 :
  (x[23:13] == 1348) ? 26'b10100111010011111011110100 :
  (x[23:13] == 1349) ? 26'b10100111001111111101111000 :
  (x[23:13] == 1350) ? 26'b10100111001100000000001000 :
  (x[23:13] == 1351) ? 26'b10100111001000000010110100 :
  (x[23:13] == 1352) ? 26'b10100111000100000101101100 :
  (x[23:13] == 1353) ? 26'b10100111000000001000110100 :
  (x[23:13] == 1354) ? 26'b10100110111100001100010000 :
  (x[23:13] == 1355) ? 26'b10100110111000010000000000 :
  (x[23:13] == 1356) ? 26'b10100110110100010100000000 :
  (x[23:13] == 1357) ? 26'b10100110110000011000010100 :
  (x[23:13] == 1358) ? 26'b10100110101100011100111000 :
  (x[23:13] == 1359) ? 26'b10100110101000100001101100 :
  (x[23:13] == 1360) ? 26'b10100110100100100110110100 :
  (x[23:13] == 1361) ? 26'b10100110100000101100001100 :
  (x[23:13] == 1362) ? 26'b10100110011100110001111000 :
  (x[23:13] == 1363) ? 26'b10100110011000110111110100 :
  (x[23:13] == 1364) ? 26'b10100110010100111110000000 :
  (x[23:13] == 1365) ? 26'b10100110010001000100100100 :
  (x[23:13] == 1366) ? 26'b10100110001101001011010100 :
  (x[23:13] == 1367) ? 26'b10100110001001010010010100 :
  (x[23:13] == 1368) ? 26'b10100110000101011001101000 :
  (x[23:13] == 1369) ? 26'b10100110000001100001010000 :
  (x[23:13] == 1370) ? 26'b10100101111101101001001000 :
  (x[23:13] == 1371) ? 26'b10100101111001110001010000 :
  (x[23:13] == 1372) ? 26'b10100101110101111001101000 :
  (x[23:13] == 1373) ? 26'b10100101110010000010010100 :
  (x[23:13] == 1374) ? 26'b10100101101110001011010000 :
  (x[23:13] == 1375) ? 26'b10100101101010010100011100 :
  (x[23:13] == 1376) ? 26'b10100101100110011101111100 :
  (x[23:13] == 1377) ? 26'b10100101100010100111101100 :
  (x[23:13] == 1378) ? 26'b10100101011110110001101100 :
  (x[23:13] == 1379) ? 26'b10100101011010111100000000 :
  (x[23:13] == 1380) ? 26'b10100101010111000110100000 :
  (x[23:13] == 1381) ? 26'b10100101010011010001010100 :
  (x[23:13] == 1382) ? 26'b10100101001111011100011000 :
  (x[23:13] == 1383) ? 26'b10100101001011100111110000 :
  (x[23:13] == 1384) ? 26'b10100101000111110011011000 :
  (x[23:13] == 1385) ? 26'b10100101000011111111010000 :
  (x[23:13] == 1386) ? 26'b10100101000000001011011000 :
  (x[23:13] == 1387) ? 26'b10100100111100010111110100 :
  (x[23:13] == 1388) ? 26'b10100100111000100100011100 :
  (x[23:13] == 1389) ? 26'b10100100110100110001011000 :
  (x[23:13] == 1390) ? 26'b10100100110000111110101000 :
  (x[23:13] == 1391) ? 26'b10100100101101001100000100 :
  (x[23:13] == 1392) ? 26'b10100100101001011001110000 :
  (x[23:13] == 1393) ? 26'b10100100100101100111110000 :
  (x[23:13] == 1394) ? 26'b10100100100001110110000000 :
  (x[23:13] == 1395) ? 26'b10100100011110000100100000 :
  (x[23:13] == 1396) ? 26'b10100100011010010011010000 :
  (x[23:13] == 1397) ? 26'b10100100010110100010010000 :
  (x[23:13] == 1398) ? 26'b10100100010010110001100100 :
  (x[23:13] == 1399) ? 26'b10100100001111000001001000 :
  (x[23:13] == 1400) ? 26'b10100100001011010000111000 :
  (x[23:13] == 1401) ? 26'b10100100000111100000111000 :
  (x[23:13] == 1402) ? 26'b10100100000011110001010000 :
  (x[23:13] == 1403) ? 26'b10100100000000000001110100 :
  (x[23:13] == 1404) ? 26'b10100011111100010010101000 :
  (x[23:13] == 1405) ? 26'b10100011111000100011101100 :
  (x[23:13] == 1406) ? 26'b10100011110100110101000000 :
  (x[23:13] == 1407) ? 26'b10100011110001000110100100 :
  (x[23:13] == 1408) ? 26'b10100011101101011000011000 :
  (x[23:13] == 1409) ? 26'b10100011101001101010100000 :
  (x[23:13] == 1410) ? 26'b10100011100101111100111000 :
  (x[23:13] == 1411) ? 26'b10100011100010001111011100 :
  (x[23:13] == 1412) ? 26'b10100011011110100010010100 :
  (x[23:13] == 1413) ? 26'b10100011011010110101011000 :
  (x[23:13] == 1414) ? 26'b10100011010111001000110000 :
  (x[23:13] == 1415) ? 26'b10100011010011011100010100 :
  (x[23:13] == 1416) ? 26'b10100011001111110000001100 :
  (x[23:13] == 1417) ? 26'b10100011001100000100010100 :
  (x[23:13] == 1418) ? 26'b10100011001000011000101000 :
  (x[23:13] == 1419) ? 26'b10100011000100101101010000 :
  (x[23:13] == 1420) ? 26'b10100011000001000010000100 :
  (x[23:13] == 1421) ? 26'b10100010111101010111001100 :
  (x[23:13] == 1422) ? 26'b10100010111001101100100000 :
  (x[23:13] == 1423) ? 26'b10100010110110000010001000 :
  (x[23:13] == 1424) ? 26'b10100010110010011000000000 :
  (x[23:13] == 1425) ? 26'b10100010101110101110000000 :
  (x[23:13] == 1426) ? 26'b10100010101011000100011000 :
  (x[23:13] == 1427) ? 26'b10100010100111011010111100 :
  (x[23:13] == 1428) ? 26'b10100010100011110001110000 :
  (x[23:13] == 1429) ? 26'b10100010100000001000110100 :
  (x[23:13] == 1430) ? 26'b10100010011100100000001000 :
  (x[23:13] == 1431) ? 26'b10100010011000110111101100 :
  (x[23:13] == 1432) ? 26'b10100010010101001111100000 :
  (x[23:13] == 1433) ? 26'b10100010010001100111100000 :
  (x[23:13] == 1434) ? 26'b10100010001101111111110100 :
  (x[23:13] == 1435) ? 26'b10100010001010011000011000 :
  (x[23:13] == 1436) ? 26'b10100010000110110001001000 :
  (x[23:13] == 1437) ? 26'b10100010000011001010001000 :
  (x[23:13] == 1438) ? 26'b10100001111111100011011000 :
  (x[23:13] == 1439) ? 26'b10100001111011111100111000 :
  (x[23:13] == 1440) ? 26'b10100001111000010110100100 :
  (x[23:13] == 1441) ? 26'b10100001110100110000100100 :
  (x[23:13] == 1442) ? 26'b10100001110001001010110000 :
  (x[23:13] == 1443) ? 26'b10100001101101100101010000 :
  (x[23:13] == 1444) ? 26'b10100001101001111111111100 :
  (x[23:13] == 1445) ? 26'b10100001100110011010111000 :
  (x[23:13] == 1446) ? 26'b10100001100010110110000000 :
  (x[23:13] == 1447) ? 26'b10100001011111010001011000 :
  (x[23:13] == 1448) ? 26'b10100001011011101101000000 :
  (x[23:13] == 1449) ? 26'b10100001011000001000111000 :
  (x[23:13] == 1450) ? 26'b10100001010100100101000000 :
  (x[23:13] == 1451) ? 26'b10100001010001000001011000 :
  (x[23:13] == 1452) ? 26'b10100001001101011101111000 :
  (x[23:13] == 1453) ? 26'b10100001001001111010110000 :
  (x[23:13] == 1454) ? 26'b10100001000110010111110000 :
  (x[23:13] == 1455) ? 26'b10100001000010110101000100 :
  (x[23:13] == 1456) ? 26'b10100000111111010010101000 :
  (x[23:13] == 1457) ? 26'b10100000111011110000010100 :
  (x[23:13] == 1458) ? 26'b10100000111000001110010100 :
  (x[23:13] == 1459) ? 26'b10100000110100101100100000 :
  (x[23:13] == 1460) ? 26'b10100000110001001011000000 :
  (x[23:13] == 1461) ? 26'b10100000101101101001101000 :
  (x[23:13] == 1462) ? 26'b10100000101010001000100100 :
  (x[23:13] == 1463) ? 26'b10100000100110100111101100 :
  (x[23:13] == 1464) ? 26'b10100000100011000111000100 :
  (x[23:13] == 1465) ? 26'b10100000011111100110101000 :
  (x[23:13] == 1466) ? 26'b10100000011100000110100000 :
  (x[23:13] == 1467) ? 26'b10100000011000100110100100 :
  (x[23:13] == 1468) ? 26'b10100000010101000110110100 :
  (x[23:13] == 1469) ? 26'b10100000010001100111010100 :
  (x[23:13] == 1470) ? 26'b10100000001110001000001000 :
  (x[23:13] == 1471) ? 26'b10100000001010101001000100 :
  (x[23:13] == 1472) ? 26'b10100000000111001010010000 :
  (x[23:13] == 1473) ? 26'b10100000000011101011101100 :
  (x[23:13] == 1474) ? 26'b10100000000000001101011000 :
  (x[23:13] == 1475) ? 26'b10011111111100101111001100 :
  (x[23:13] == 1476) ? 26'b10011111111001010001010100 :
  (x[23:13] == 1477) ? 26'b10011111110101110011101000 :
  (x[23:13] == 1478) ? 26'b10011111110010010110001100 :
  (x[23:13] == 1479) ? 26'b10011111101110111001000000 :
  (x[23:13] == 1480) ? 26'b10011111101011011100000000 :
  (x[23:13] == 1481) ? 26'b10011111100111111111001100 :
  (x[23:13] == 1482) ? 26'b10011111100100100010101000 :
  (x[23:13] == 1483) ? 26'b10011111100001000110010100 :
  (x[23:13] == 1484) ? 26'b10011111011101101010001100 :
  (x[23:13] == 1485) ? 26'b10011111011010001110010100 :
  (x[23:13] == 1486) ? 26'b10011111010110110010101000 :
  (x[23:13] == 1487) ? 26'b10011111010011010111010000 :
  (x[23:13] == 1488) ? 26'b10011111001111111100000000 :
  (x[23:13] == 1489) ? 26'b10011111001100100001000000 :
  (x[23:13] == 1490) ? 26'b10011111001001000110010000 :
  (x[23:13] == 1491) ? 26'b10011111000101101011101100 :
  (x[23:13] == 1492) ? 26'b10011111000010010001011000 :
  (x[23:13] == 1493) ? 26'b10011110111110110111010000 :
  (x[23:13] == 1494) ? 26'b10011110111011011101010100 :
  (x[23:13] == 1495) ? 26'b10011110111000000011101000 :
  (x[23:13] == 1496) ? 26'b10011110110100101010001100 :
  (x[23:13] == 1497) ? 26'b10011110110001010000111100 :
  (x[23:13] == 1498) ? 26'b10011110101101110111111100 :
  (x[23:13] == 1499) ? 26'b10011110101010011111001000 :
  (x[23:13] == 1500) ? 26'b10011110100111000110100000 :
  (x[23:13] == 1501) ? 26'b10011110100011101110001000 :
  (x[23:13] == 1502) ? 26'b10011110100000010110000000 :
  (x[23:13] == 1503) ? 26'b10011110011100111110000000 :
  (x[23:13] == 1504) ? 26'b10011110011001100110010100 :
  (x[23:13] == 1505) ? 26'b10011110010110001110110000 :
  (x[23:13] == 1506) ? 26'b10011110010010110111100000 :
  (x[23:13] == 1507) ? 26'b10011110001111100000011000 :
  (x[23:13] == 1508) ? 26'b10011110001100001001100000 :
  (x[23:13] == 1509) ? 26'b10011110001000110010111000 :
  (x[23:13] == 1510) ? 26'b10011110000101011100011100 :
  (x[23:13] == 1511) ? 26'b10011110000010000110001100 :
  (x[23:13] == 1512) ? 26'b10011101111110110000001100 :
  (x[23:13] == 1513) ? 26'b10011101111011011010011000 :
  (x[23:13] == 1514) ? 26'b10011101111000000100110000 :
  (x[23:13] == 1515) ? 26'b10011101110100101111011000 :
  (x[23:13] == 1516) ? 26'b10011101110001011010010000 :
  (x[23:13] == 1517) ? 26'b10011101101110000101010000 :
  (x[23:13] == 1518) ? 26'b10011101101010110000100000 :
  (x[23:13] == 1519) ? 26'b10011101100111011100000000 :
  (x[23:13] == 1520) ? 26'b10011101100100000111101000 :
  (x[23:13] == 1521) ? 26'b10011101100000110011100000 :
  (x[23:13] == 1522) ? 26'b10011101011101011111101000 :
  (x[23:13] == 1523) ? 26'b10011101011010001011111000 :
  (x[23:13] == 1524) ? 26'b10011101010110111000011000 :
  (x[23:13] == 1525) ? 26'b10011101010011100101001000 :
  (x[23:13] == 1526) ? 26'b10011101010000010010000000 :
  (x[23:13] == 1527) ? 26'b10011101001100111111001000 :
  (x[23:13] == 1528) ? 26'b10011101001001101100100000 :
  (x[23:13] == 1529) ? 26'b10011101000110011010000000 :
  (x[23:13] == 1530) ? 26'b10011101000011000111110000 :
  (x[23:13] == 1531) ? 26'b10011100111111110101110000 :
  (x[23:13] == 1532) ? 26'b10011100111100100011111000 :
  (x[23:13] == 1533) ? 26'b10011100111001010010010000 :
  (x[23:13] == 1534) ? 26'b10011100110110000000110100 :
  (x[23:13] == 1535) ? 26'b10011100110010101111101000 :
  (x[23:13] == 1536) ? 26'b10011100101111011110100000 :
  (x[23:13] == 1537) ? 26'b10011100101100001101110000 :
  (x[23:13] == 1538) ? 26'b10011100101000111101001000 :
  (x[23:13] == 1539) ? 26'b10011100100101101100101100 :
  (x[23:13] == 1540) ? 26'b10011100100010011100100000 :
  (x[23:13] == 1541) ? 26'b10011100011111001100100000 :
  (x[23:13] == 1542) ? 26'b10011100011011111100101100 :
  (x[23:13] == 1543) ? 26'b10011100011000101101001000 :
  (x[23:13] == 1544) ? 26'b10011100010101011101101100 :
  (x[23:13] == 1545) ? 26'b10011100010010001110100000 :
  (x[23:13] == 1546) ? 26'b10011100001110111111100000 :
  (x[23:13] == 1547) ? 26'b10011100001011110000101100 :
  (x[23:13] == 1548) ? 26'b10011100001000100010001000 :
  (x[23:13] == 1549) ? 26'b10011100000101010011101100 :
  (x[23:13] == 1550) ? 26'b10011100000010000101100000 :
  (x[23:13] == 1551) ? 26'b10011011111110110111100000 :
  (x[23:13] == 1552) ? 26'b10011011111011101001101100 :
  (x[23:13] == 1553) ? 26'b10011011111000011100001000 :
  (x[23:13] == 1554) ? 26'b10011011110101001110101100 :
  (x[23:13] == 1555) ? 26'b10011011110010000001100000 :
  (x[23:13] == 1556) ? 26'b10011011101110110100100000 :
  (x[23:13] == 1557) ? 26'b10011011101011100111101000 :
  (x[23:13] == 1558) ? 26'b10011011101000011011000100 :
  (x[23:13] == 1559) ? 26'b10011011100101001110101100 :
  (x[23:13] == 1560) ? 26'b10011011100010000010011100 :
  (x[23:13] == 1561) ? 26'b10011011011110110110011000 :
  (x[23:13] == 1562) ? 26'b10011011011011101010100100 :
  (x[23:13] == 1563) ? 26'b10011011011000011110111100 :
  (x[23:13] == 1564) ? 26'b10011011010101010011100000 :
  (x[23:13] == 1565) ? 26'b10011011010010001000010000 :
  (x[23:13] == 1566) ? 26'b10011011001110111101010000 :
  (x[23:13] == 1567) ? 26'b10011011001011110010011000 :
  (x[23:13] == 1568) ? 26'b10011011001000100111110000 :
  (x[23:13] == 1569) ? 26'b10011011000101011101010000 :
  (x[23:13] == 1570) ? 26'b10011011000010010011000000 :
  (x[23:13] == 1571) ? 26'b10011010111111001000111000 :
  (x[23:13] == 1572) ? 26'b10011010111011111111000100 :
  (x[23:13] == 1573) ? 26'b10011010111000110101011000 :
  (x[23:13] == 1574) ? 26'b10011010110101101011110100 :
  (x[23:13] == 1575) ? 26'b10011010110010100010100100 :
  (x[23:13] == 1576) ? 26'b10011010101111011001011000 :
  (x[23:13] == 1577) ? 26'b10011010101100010000100000 :
  (x[23:13] == 1578) ? 26'b10011010101001000111110000 :
  (x[23:13] == 1579) ? 26'b10011010100101111111001100 :
  (x[23:13] == 1580) ? 26'b10011010100010110110111000 :
  (x[23:13] == 1581) ? 26'b10011010011111101110101100 :
  (x[23:13] == 1582) ? 26'b10011010011100100110110000 :
  (x[23:13] == 1583) ? 26'b10011010011001011110111100 :
  (x[23:13] == 1584) ? 26'b10011010010110010111011000 :
  (x[23:13] == 1585) ? 26'b10011010010011001111111100 :
  (x[23:13] == 1586) ? 26'b10011010010000001000110000 :
  (x[23:13] == 1587) ? 26'b10011010001101000001101100 :
  (x[23:13] == 1588) ? 26'b10011010001001111010111000 :
  (x[23:13] == 1589) ? 26'b10011010000110110100001100 :
  (x[23:13] == 1590) ? 26'b10011010000011101101110000 :
  (x[23:13] == 1591) ? 26'b10011010000000100111011100 :
  (x[23:13] == 1592) ? 26'b10011001111101100001011000 :
  (x[23:13] == 1593) ? 26'b10011001111010011011011100 :
  (x[23:13] == 1594) ? 26'b10011001110111010101110000 :
  (x[23:13] == 1595) ? 26'b10011001110100010000001100 :
  (x[23:13] == 1596) ? 26'b10011001110001001010111000 :
  (x[23:13] == 1597) ? 26'b10011001101110000101101100 :
  (x[23:13] == 1598) ? 26'b10011001101011000000110000 :
  (x[23:13] == 1599) ? 26'b10011001100111111011111000 :
  (x[23:13] == 1600) ? 26'b10011001100100110111010100 :
  (x[23:13] == 1601) ? 26'b10011001100001110010111000 :
  (x[23:13] == 1602) ? 26'b10011001011110101110101000 :
  (x[23:13] == 1603) ? 26'b10011001011011101010101000 :
  (x[23:13] == 1604) ? 26'b10011001011000100110110000 :
  (x[23:13] == 1605) ? 26'b10011001010101100011000000 :
  (x[23:13] == 1606) ? 26'b10011001010010011111100100 :
  (x[23:13] == 1607) ? 26'b10011001001111011100010000 :
  (x[23:13] == 1608) ? 26'b10011001001100011001000100 :
  (x[23:13] == 1609) ? 26'b10011001001001010110000100 :
  (x[23:13] == 1610) ? 26'b10011001000110010011010100 :
  (x[23:13] == 1611) ? 26'b10011001000011010000110000 :
  (x[23:13] == 1612) ? 26'b10011001000000001110010100 :
  (x[23:13] == 1613) ? 26'b10011000111101001100001000 :
  (x[23:13] == 1614) ? 26'b10011000111010001010000000 :
  (x[23:13] == 1615) ? 26'b10011000110111001000001000 :
  (x[23:13] == 1616) ? 26'b10011000110100000110011100 :
  (x[23:13] == 1617) ? 26'b10011000110001000100111100 :
  (x[23:13] == 1618) ? 26'b10011000101110000011101000 :
  (x[23:13] == 1619) ? 26'b10011000101011000010011100 :
  (x[23:13] == 1620) ? 26'b10011000101000000001011100 :
  (x[23:13] == 1621) ? 26'b10011000100101000000101000 :
  (x[23:13] == 1622) ? 26'b10011000100010000000000100 :
  (x[23:13] == 1623) ? 26'b10011000011110111111100100 :
  (x[23:13] == 1624) ? 26'b10011000011011111111011000 :
  (x[23:13] == 1625) ? 26'b10011000011000111111010000 :
  (x[23:13] == 1626) ? 26'b10011000010101111111011000 :
  (x[23:13] == 1627) ? 26'b10011000010010111111100100 :
  (x[23:13] == 1628) ? 26'b10011000010000000000000100 :
  (x[23:13] == 1629) ? 26'b10011000001101000000101000 :
  (x[23:13] == 1630) ? 26'b10011000001010000001011100 :
  (x[23:13] == 1631) ? 26'b10011000000111000010011100 :
  (x[23:13] == 1632) ? 26'b10011000000100000011100100 :
  (x[23:13] == 1633) ? 26'b10011000000001000100111000 :
  (x[23:13] == 1634) ? 26'b10010111111110000110011000 :
  (x[23:13] == 1635) ? 26'b10010111111011001000000100 :
  (x[23:13] == 1636) ? 26'b10010111111000001001111000 :
  (x[23:13] == 1637) ? 26'b10010111110101001011111000 :
  (x[23:13] == 1638) ? 26'b10010111110010001110001000 :
  (x[23:13] == 1639) ? 26'b10010111101111010000100000 :
  (x[23:13] == 1640) ? 26'b10010111101100010011000000 :
  (x[23:13] == 1641) ? 26'b10010111101001010101110000 :
  (x[23:13] == 1642) ? 26'b10010111100110011000101000 :
  (x[23:13] == 1643) ? 26'b10010111100011011011101100 :
  (x[23:13] == 1644) ? 26'b10010111100000011110111100 :
  (x[23:13] == 1645) ? 26'b10010111011101100010010100 :
  (x[23:13] == 1646) ? 26'b10010111011010100101111000 :
  (x[23:13] == 1647) ? 26'b10010111010111101001101000 :
  (x[23:13] == 1648) ? 26'b10010111010100101101100100 :
  (x[23:13] == 1649) ? 26'b10010111010001110001101000 :
  (x[23:13] == 1650) ? 26'b10010111001110110101111000 :
  (x[23:13] == 1651) ? 26'b10010111001011111010011000 :
  (x[23:13] == 1652) ? 26'b10010111001000111110111100 :
  (x[23:13] == 1653) ? 26'b10010111000110000011110000 :
  (x[23:13] == 1654) ? 26'b10010111000011001000101000 :
  (x[23:13] == 1655) ? 26'b10010111000000001101110000 :
  (x[23:13] == 1656) ? 26'b10010110111101010011000100 :
  (x[23:13] == 1657) ? 26'b10010110111010011000100000 :
  (x[23:13] == 1658) ? 26'b10010110110111011110001000 :
  (x[23:13] == 1659) ? 26'b10010110110100100011111000 :
  (x[23:13] == 1660) ? 26'b10010110110001101001111000 :
  (x[23:13] == 1661) ? 26'b10010110101110110000000000 :
  (x[23:13] == 1662) ? 26'b10010110101011110110010000 :
  (x[23:13] == 1663) ? 26'b10010110101000111100110000 :
  (x[23:13] == 1664) ? 26'b10010110100110000011011000 :
  (x[23:13] == 1665) ? 26'b10010110100011001010001000 :
  (x[23:13] == 1666) ? 26'b10010110100000010001001000 :
  (x[23:13] == 1667) ? 26'b10010110011101011000010000 :
  (x[23:13] == 1668) ? 26'b10010110011010011111100000 :
  (x[23:13] == 1669) ? 26'b10010110010111100111000000 :
  (x[23:13] == 1670) ? 26'b10010110010100101110101000 :
  (x[23:13] == 1671) ? 26'b10010110010001110110011000 :
  (x[23:13] == 1672) ? 26'b10010110001110111110011000 :
  (x[23:13] == 1673) ? 26'b10010110001100000110100000 :
  (x[23:13] == 1674) ? 26'b10010110001001001110110000 :
  (x[23:13] == 1675) ? 26'b10010110000110010111001100 :
  (x[23:13] == 1676) ? 26'b10010110000011011111110000 :
  (x[23:13] == 1677) ? 26'b10010110000000101000101000 :
  (x[23:13] == 1678) ? 26'b10010101111101110001100000 :
  (x[23:13] == 1679) ? 26'b10010101111010111010101000 :
  (x[23:13] == 1680) ? 26'b10010101111000000011111000 :
  (x[23:13] == 1681) ? 26'b10010101110101001101011000 :
  (x[23:13] == 1682) ? 26'b10010101110010010110111000 :
  (x[23:13] == 1683) ? 26'b10010101101111100000101000 :
  (x[23:13] == 1684) ? 26'b10010101101100101010101000 :
  (x[23:13] == 1685) ? 26'b10010101101001110100101100 :
  (x[23:13] == 1686) ? 26'b10010101100110111110111000 :
  (x[23:13] == 1687) ? 26'b10010101100100001001010100 :
  (x[23:13] == 1688) ? 26'b10010101100001010011111000 :
  (x[23:13] == 1689) ? 26'b10010101011110011110100100 :
  (x[23:13] == 1690) ? 26'b10010101011011101001100000 :
  (x[23:13] == 1691) ? 26'b10010101011000110100100000 :
  (x[23:13] == 1692) ? 26'b10010101010101111111110000 :
  (x[23:13] == 1693) ? 26'b10010101010011001011001000 :
  (x[23:13] == 1694) ? 26'b10010101010000010110101000 :
  (x[23:13] == 1695) ? 26'b10010101001101100010010100 :
  (x[23:13] == 1696) ? 26'b10010101001010101110001100 :
  (x[23:13] == 1697) ? 26'b10010101000111111010001100 :
  (x[23:13] == 1698) ? 26'b10010101000101000110011000 :
  (x[23:13] == 1699) ? 26'b10010101000010010010101100 :
  (x[23:13] == 1700) ? 26'b10010100111111011111001000 :
  (x[23:13] == 1701) ? 26'b10010100111100101011110000 :
  (x[23:13] == 1702) ? 26'b10010100111001111000100100 :
  (x[23:13] == 1703) ? 26'b10010100110111000101100100 :
  (x[23:13] == 1704) ? 26'b10010100110100010010101100 :
  (x[23:13] == 1705) ? 26'b10010100110001011111111100 :
  (x[23:13] == 1706) ? 26'b10010100101110101101011000 :
  (x[23:13] == 1707) ? 26'b10010100101011111010111100 :
  (x[23:13] == 1708) ? 26'b10010100101001001000101100 :
  (x[23:13] == 1709) ? 26'b10010100100110010110101000 :
  (x[23:13] == 1710) ? 26'b10010100100011100100101000 :
  (x[23:13] == 1711) ? 26'b10010100100000110010111000 :
  (x[23:13] == 1712) ? 26'b10010100011110000001001100 :
  (x[23:13] == 1713) ? 26'b10010100011011001111110000 :
  (x[23:13] == 1714) ? 26'b10010100011000011110011000 :
  (x[23:13] == 1715) ? 26'b10010100010101101101010000 :
  (x[23:13] == 1716) ? 26'b10010100010010111100010000 :
  (x[23:13] == 1717) ? 26'b10010100010000001011011000 :
  (x[23:13] == 1718) ? 26'b10010100001101011010101100 :
  (x[23:13] == 1719) ? 26'b10010100001010101010001000 :
  (x[23:13] == 1720) ? 26'b10010100000111111001110000 :
  (x[23:13] == 1721) ? 26'b10010100000101001001100000 :
  (x[23:13] == 1722) ? 26'b10010100000010011001011000 :
  (x[23:13] == 1723) ? 26'b10010011111111101001011100 :
  (x[23:13] == 1724) ? 26'b10010011111100111001101000 :
  (x[23:13] == 1725) ? 26'b10010011111010001010000100 :
  (x[23:13] == 1726) ? 26'b10010011110111011010100100 :
  (x[23:13] == 1727) ? 26'b10010011110100101011010000 :
  (x[23:13] == 1728) ? 26'b10010011110001111100000100 :
  (x[23:13] == 1729) ? 26'b10010011101111001101000100 :
  (x[23:13] == 1730) ? 26'b10010011101100011110001000 :
  (x[23:13] == 1731) ? 26'b10010011101001101111011100 :
  (x[23:13] == 1732) ? 26'b10010011100111000000111000 :
  (x[23:13] == 1733) ? 26'b10010011100100010010100000 :
  (x[23:13] == 1734) ? 26'b10010011100001100100010000 :
  (x[23:13] == 1735) ? 26'b10010011011110110110001000 :
  (x[23:13] == 1736) ? 26'b10010011011100001000001000 :
  (x[23:13] == 1737) ? 26'b10010011011001011010010100 :
  (x[23:13] == 1738) ? 26'b10010011010110101100101000 :
  (x[23:13] == 1739) ? 26'b10010011010011111111001100 :
  (x[23:13] == 1740) ? 26'b10010011010001010001110000 :
  (x[23:13] == 1741) ? 26'b10010011001110100100100100 :
  (x[23:13] == 1742) ? 26'b10010011001011110111100000 :
  (x[23:13] == 1743) ? 26'b10010011001001001010101000 :
  (x[23:13] == 1744) ? 26'b10010011000110011101110100 :
  (x[23:13] == 1745) ? 26'b10010011000011110001010000 :
  (x[23:13] == 1746) ? 26'b10010011000001000100110000 :
  (x[23:13] == 1747) ? 26'b10010010111110011000011000 :
  (x[23:13] == 1748) ? 26'b10010010111011101100010000 :
  (x[23:13] == 1749) ? 26'b10010010111001000000001100 :
  (x[23:13] == 1750) ? 26'b10010010110110010100010100 :
  (x[23:13] == 1751) ? 26'b10010010110011101000101000 :
  (x[23:13] == 1752) ? 26'b10010010110000111101000000 :
  (x[23:13] == 1753) ? 26'b10010010101110010001100100 :
  (x[23:13] == 1754) ? 26'b10010010101011100110010100 :
  (x[23:13] == 1755) ? 26'b10010010101000111011001000 :
  (x[23:13] == 1756) ? 26'b10010010100110010000001000 :
  (x[23:13] == 1757) ? 26'b10010010100011100101010100 :
  (x[23:13] == 1758) ? 26'b10010010100000111010100100 :
  (x[23:13] == 1759) ? 26'b10010010011110010000000000 :
  (x[23:13] == 1760) ? 26'b10010010011011100101101000 :
  (x[23:13] == 1761) ? 26'b10010010011000111011010100 :
  (x[23:13] == 1762) ? 26'b10010010010110010001001100 :
  (x[23:13] == 1763) ? 26'b10010010010011100111010000 :
  (x[23:13] == 1764) ? 26'b10010010010000111101011000 :
  (x[23:13] == 1765) ? 26'b10010010001110010011101100 :
  (x[23:13] == 1766) ? 26'b10010010001011101010001000 :
  (x[23:13] == 1767) ? 26'b10010010001001000000110000 :
  (x[23:13] == 1768) ? 26'b10010010000110010111100000 :
  (x[23:13] == 1769) ? 26'b10010010000011101110011000 :
  (x[23:13] == 1770) ? 26'b10010010000001000101011000 :
  (x[23:13] == 1771) ? 26'b10010001111110011100100100 :
  (x[23:13] == 1772) ? 26'b10010001111011110011111000 :
  (x[23:13] == 1773) ? 26'b10010001111001001011010100 :
  (x[23:13] == 1774) ? 26'b10010001110110100010111000 :
  (x[23:13] == 1775) ? 26'b10010001110011111010101100 :
  (x[23:13] == 1776) ? 26'b10010001110001010010100000 :
  (x[23:13] == 1777) ? 26'b10010001101110101010100100 :
  (x[23:13] == 1778) ? 26'b10010001101100000010110000 :
  (x[23:13] == 1779) ? 26'b10010001101001011011000100 :
  (x[23:13] == 1780) ? 26'b10010001100110110011100000 :
  (x[23:13] == 1781) ? 26'b10010001100100001100000100 :
  (x[23:13] == 1782) ? 26'b10010001100001100100110000 :
  (x[23:13] == 1783) ? 26'b10010001011110111101101100 :
  (x[23:13] == 1784) ? 26'b10010001011100010110101000 :
  (x[23:13] == 1785) ? 26'b10010001011001101111110100 :
  (x[23:13] == 1786) ? 26'b10010001010111001001001000 :
  (x[23:13] == 1787) ? 26'b10010001010100100010100100 :
  (x[23:13] == 1788) ? 26'b10010001010001111100001000 :
  (x[23:13] == 1789) ? 26'b10010001001111010101110100 :
  (x[23:13] == 1790) ? 26'b10010001001100101111101000 :
  (x[23:13] == 1791) ? 26'b10010001001010001001101100 :
  (x[23:13] == 1792) ? 26'b10010001000111100011110000 :
  (x[23:13] == 1793) ? 26'b10010001000100111110000100 :
  (x[23:13] == 1794) ? 26'b10010001000010011000100000 :
  (x[23:13] == 1795) ? 26'b10010000111111110011000000 :
  (x[23:13] == 1796) ? 26'b10010000111101001101101100 :
  (x[23:13] == 1797) ? 26'b10010000111010101000100000 :
  (x[23:13] == 1798) ? 26'b10010000111000000011100000 :
  (x[23:13] == 1799) ? 26'b10010000110101011110100100 :
  (x[23:13] == 1800) ? 26'b10010000110010111001110100 :
  (x[23:13] == 1801) ? 26'b10010000110000010101001000 :
  (x[23:13] == 1802) ? 26'b10010000101101110000101000 :
  (x[23:13] == 1803) ? 26'b10010000101011001100010100 :
  (x[23:13] == 1804) ? 26'b10010000101000101000001000 :
  (x[23:13] == 1805) ? 26'b10010000100110000100000000 :
  (x[23:13] == 1806) ? 26'b10010000100011100000000100 :
  (x[23:13] == 1807) ? 26'b10010000100000111100010000 :
  (x[23:13] == 1808) ? 26'b10010000011110011000100100 :
  (x[23:13] == 1809) ? 26'b10010000011011110101000000 :
  (x[23:13] == 1810) ? 26'b10010000011001010001101000 :
  (x[23:13] == 1811) ? 26'b10010000010110101110011000 :
  (x[23:13] == 1812) ? 26'b10010000010100001011010000 :
  (x[23:13] == 1813) ? 26'b10010000010001101000010000 :
  (x[23:13] == 1814) ? 26'b10010000001111000101011000 :
  (x[23:13] == 1815) ? 26'b10010000001100100010101000 :
  (x[23:13] == 1816) ? 26'b10010000001010000000000000 :
  (x[23:13] == 1817) ? 26'b10010000000111011101100100 :
  (x[23:13] == 1818) ? 26'b10010000000100111011010000 :
  (x[23:13] == 1819) ? 26'b10010000000010011001000100 :
  (x[23:13] == 1820) ? 26'b10001111111111110111000000 :
  (x[23:13] == 1821) ? 26'b10001111111101010101001000 :
  (x[23:13] == 1822) ? 26'b10001111111010110011010000 :
  (x[23:13] == 1823) ? 26'b10001111111000010001101000 :
  (x[23:13] == 1824) ? 26'b10001111110101110000000100 :
  (x[23:13] == 1825) ? 26'b10001111110011001110101100 :
  (x[23:13] == 1826) ? 26'b10001111110000101101011100 :
  (x[23:13] == 1827) ? 26'b10001111101110001100010100 :
  (x[23:13] == 1828) ? 26'b10001111101011101011010100 :
  (x[23:13] == 1829) ? 26'b10001111101001001010011100 :
  (x[23:13] == 1830) ? 26'b10001111100110101001101100 :
  (x[23:13] == 1831) ? 26'b10001111100100001001001000 :
  (x[23:13] == 1832) ? 26'b10001111100001101000101000 :
  (x[23:13] == 1833) ? 26'b10001111011111001000010100 :
  (x[23:13] == 1834) ? 26'b10001111011100101000000100 :
  (x[23:13] == 1835) ? 26'b10001111011010001000000100 :
  (x[23:13] == 1836) ? 26'b10001111010111101000000100 :
  (x[23:13] == 1837) ? 26'b10001111010101001000010000 :
  (x[23:13] == 1838) ? 26'b10001111010010101000100100 :
  (x[23:13] == 1839) ? 26'b10001111010000001001000100 :
  (x[23:13] == 1840) ? 26'b10001111001101101001100100 :
  (x[23:13] == 1841) ? 26'b10001111001011001010010100 :
  (x[23:13] == 1842) ? 26'b10001111001000101011001000 :
  (x[23:13] == 1843) ? 26'b10001111000110001100001000 :
  (x[23:13] == 1844) ? 26'b10001111000011101101001100 :
  (x[23:13] == 1845) ? 26'b10001111000001001110011100 :
  (x[23:13] == 1846) ? 26'b10001110111110101111110000 :
  (x[23:13] == 1847) ? 26'b10001110111100010001010000 :
  (x[23:13] == 1848) ? 26'b10001110111001110010111000 :
  (x[23:13] == 1849) ? 26'b10001110110111010100101000 :
  (x[23:13] == 1850) ? 26'b10001110110100110110100000 :
  (x[23:13] == 1851) ? 26'b10001110110010011000100000 :
  (x[23:13] == 1852) ? 26'b10001110101111111010101000 :
  (x[23:13] == 1853) ? 26'b10001110101101011100111000 :
  (x[23:13] == 1854) ? 26'b10001110101010111111010000 :
  (x[23:13] == 1855) ? 26'b10001110101000100001110000 :
  (x[23:13] == 1856) ? 26'b10001110100110000100011000 :
  (x[23:13] == 1857) ? 26'b10001110100011100111001000 :
  (x[23:13] == 1858) ? 26'b10001110100001001010000000 :
  (x[23:13] == 1859) ? 26'b10001110011110101101000000 :
  (x[23:13] == 1860) ? 26'b10001110011100010000001000 :
  (x[23:13] == 1861) ? 26'b10001110011001110011011100 :
  (x[23:13] == 1862) ? 26'b10001110010111010110110100 :
  (x[23:13] == 1863) ? 26'b10001110010100111010010100 :
  (x[23:13] == 1864) ? 26'b10001110010010011110000000 :
  (x[23:13] == 1865) ? 26'b10001110010000000001110000 :
  (x[23:13] == 1866) ? 26'b10001110001101100101101000 :
  (x[23:13] == 1867) ? 26'b10001110001011001001101000 :
  (x[23:13] == 1868) ? 26'b10001110001000101101110100 :
  (x[23:13] == 1869) ? 26'b10001110000110010010000100 :
  (x[23:13] == 1870) ? 26'b10001110000011110110100000 :
  (x[23:13] == 1871) ? 26'b10001110000001011011000000 :
  (x[23:13] == 1872) ? 26'b10001101111110111111101100 :
  (x[23:13] == 1873) ? 26'b10001101111100100100011100 :
  (x[23:13] == 1874) ? 26'b10001101111010001001010100 :
  (x[23:13] == 1875) ? 26'b10001101110111101110011000 :
  (x[23:13] == 1876) ? 26'b10001101110101010011100000 :
  (x[23:13] == 1877) ? 26'b10001101110010111000110000 :
  (x[23:13] == 1878) ? 26'b10001101110000011110001000 :
  (x[23:13] == 1879) ? 26'b10001101101110000011101000 :
  (x[23:13] == 1880) ? 26'b10001101101011101001010000 :
  (x[23:13] == 1881) ? 26'b10001101101001001111000100 :
  (x[23:13] == 1882) ? 26'b10001101100110110100111100 :
  (x[23:13] == 1883) ? 26'b10001101100100011010111100 :
  (x[23:13] == 1884) ? 26'b10001101100010000001000100 :
  (x[23:13] == 1885) ? 26'b10001101011111100111010100 :
  (x[23:13] == 1886) ? 26'b10001101011101001101101100 :
  (x[23:13] == 1887) ? 26'b10001101011010110100001100 :
  (x[23:13] == 1888) ? 26'b10001101011000011010110100 :
  (x[23:13] == 1889) ? 26'b10001101010110000001100000 :
  (x[23:13] == 1890) ? 26'b10001101010011101000011000 :
  (x[23:13] == 1891) ? 26'b10001101010001001111011000 :
  (x[23:13] == 1892) ? 26'b10001101001110110110100000 :
  (x[23:13] == 1893) ? 26'b10001101001100011101110000 :
  (x[23:13] == 1894) ? 26'b10001101001010000101000100 :
  (x[23:13] == 1895) ? 26'b10001101000111101100100000 :
  (x[23:13] == 1896) ? 26'b10001101000101010100000100 :
  (x[23:13] == 1897) ? 26'b10001101000010111011110100 :
  (x[23:13] == 1898) ? 26'b10001101000000100011101000 :
  (x[23:13] == 1899) ? 26'b10001100111110001011100100 :
  (x[23:13] == 1900) ? 26'b10001100111011110011101000 :
  (x[23:13] == 1901) ? 26'b10001100111001011011110100 :
  (x[23:13] == 1902) ? 26'b10001100110111000100001000 :
  (x[23:13] == 1903) ? 26'b10001100110100101100100100 :
  (x[23:13] == 1904) ? 26'b10001100110010010101001000 :
  (x[23:13] == 1905) ? 26'b10001100101111111101110000 :
  (x[23:13] == 1906) ? 26'b10001100101101100110100100 :
  (x[23:13] == 1907) ? 26'b10001100101011001111100000 :
  (x[23:13] == 1908) ? 26'b10001100101000111000100000 :
  (x[23:13] == 1909) ? 26'b10001100100110100001101000 :
  (x[23:13] == 1910) ? 26'b10001100100100001010111000 :
  (x[23:13] == 1911) ? 26'b10001100100001110100010000 :
  (x[23:13] == 1912) ? 26'b10001100011111011101110000 :
  (x[23:13] == 1913) ? 26'b10001100011101000111011000 :
  (x[23:13] == 1914) ? 26'b10001100011010110001001000 :
  (x[23:13] == 1915) ? 26'b10001100011000011011000000 :
  (x[23:13] == 1916) ? 26'b10001100010110000100111100 :
  (x[23:13] == 1917) ? 26'b10001100010011101111000000 :
  (x[23:13] == 1918) ? 26'b10001100010001011001001100 :
  (x[23:13] == 1919) ? 26'b10001100001111000011100000 :
  (x[23:13] == 1920) ? 26'b10001100001100101101111100 :
  (x[23:13] == 1921) ? 26'b10001100001010011000100000 :
  (x[23:13] == 1922) ? 26'b10001100001000000011001100 :
  (x[23:13] == 1923) ? 26'b10001100000101101110000000 :
  (x[23:13] == 1924) ? 26'b10001100000011011000111000 :
  (x[23:13] == 1925) ? 26'b10001100000001000011111000 :
  (x[23:13] == 1926) ? 26'b10001011111110101111000000 :
  (x[23:13] == 1927) ? 26'b10001011111100011010010000 :
  (x[23:13] == 1928) ? 26'b10001011111010000101101000 :
  (x[23:13] == 1929) ? 26'b10001011110111110001001000 :
  (x[23:13] == 1930) ? 26'b10001011110101011100101100 :
  (x[23:13] == 1931) ? 26'b10001011110011001000011100 :
  (x[23:13] == 1932) ? 26'b10001011110000110100010000 :
  (x[23:13] == 1933) ? 26'b10001011101110100000001100 :
  (x[23:13] == 1934) ? 26'b10001011101100001100010000 :
  (x[23:13] == 1935) ? 26'b10001011101001111000011100 :
  (x[23:13] == 1936) ? 26'b10001011100111100100101100 :
  (x[23:13] == 1937) ? 26'b10001011100101010001001000 :
  (x[23:13] == 1938) ? 26'b10001011100010111101101000 :
  (x[23:13] == 1939) ? 26'b10001011100000101010010000 :
  (x[23:13] == 1940) ? 26'b10001011011110010111000000 :
  (x[23:13] == 1941) ? 26'b10001011011100000011111000 :
  (x[23:13] == 1942) ? 26'b10001011011001110000110100 :
  (x[23:13] == 1943) ? 26'b10001011010111011101111000 :
  (x[23:13] == 1944) ? 26'b10001011010101001011001000 :
  (x[23:13] == 1945) ? 26'b10001011010010111000011100 :
  (x[23:13] == 1946) ? 26'b10001011010000100101111000 :
  (x[23:13] == 1947) ? 26'b10001011001110010011011000 :
  (x[23:13] == 1948) ? 26'b10001011001100000001000000 :
  (x[23:13] == 1949) ? 26'b10001011001001101110110000 :
  (x[23:13] == 1950) ? 26'b10001011000111011100101000 :
  (x[23:13] == 1951) ? 26'b10001011000101001010101000 :
  (x[23:13] == 1952) ? 26'b10001011000010111000110000 :
  (x[23:13] == 1953) ? 26'b10001011000000100110111100 :
  (x[23:13] == 1954) ? 26'b10001010111110010101010000 :
  (x[23:13] == 1955) ? 26'b10001010111100000011101100 :
  (x[23:13] == 1956) ? 26'b10001010111001110010010000 :
  (x[23:13] == 1957) ? 26'b10001010110111100000111000 :
  (x[23:13] == 1958) ? 26'b10001010110101001111101100 :
  (x[23:13] == 1959) ? 26'b10001010110010111110100100 :
  (x[23:13] == 1960) ? 26'b10001010110000101101100000 :
  (x[23:13] == 1961) ? 26'b10001010101110011100101000 :
  (x[23:13] == 1962) ? 26'b10001010101100001011110100 :
  (x[23:13] == 1963) ? 26'b10001010101001111011001100 :
  (x[23:13] == 1964) ? 26'b10001010100111101010101000 :
  (x[23:13] == 1965) ? 26'b10001010100101011010001000 :
  (x[23:13] == 1966) ? 26'b10001010100011001001110100 :
  (x[23:13] == 1967) ? 26'b10001010100000111001100100 :
  (x[23:13] == 1968) ? 26'b10001010011110101001011100 :
  (x[23:13] == 1969) ? 26'b10001010011100011001011100 :
  (x[23:13] == 1970) ? 26'b10001010011010001001100000 :
  (x[23:13] == 1971) ? 26'b10001010010111111001110000 :
  (x[23:13] == 1972) ? 26'b10001010010101101010000100 :
  (x[23:13] == 1973) ? 26'b10001010010011011010100000 :
  (x[23:13] == 1974) ? 26'b10001010010001001011000000 :
  (x[23:13] == 1975) ? 26'b10001010001110111011101000 :
  (x[23:13] == 1976) ? 26'b10001010001100101100011000 :
  (x[23:13] == 1977) ? 26'b10001010001010011101010000 :
  (x[23:13] == 1978) ? 26'b10001010001000001110001100 :
  (x[23:13] == 1979) ? 26'b10001010000101111111010000 :
  (x[23:13] == 1980) ? 26'b10001010000011110000011100 :
  (x[23:13] == 1981) ? 26'b10001010000001100001110000 :
  (x[23:13] == 1982) ? 26'b10001001111111010011001000 :
  (x[23:13] == 1983) ? 26'b10001001111101000100101000 :
  (x[23:13] == 1984) ? 26'b10001001111010110110010000 :
  (x[23:13] == 1985) ? 26'b10001001111000101000000000 :
  (x[23:13] == 1986) ? 26'b10001001110110011001110100 :
  (x[23:13] == 1987) ? 26'b10001001110100001011110000 :
  (x[23:13] == 1988) ? 26'b10001001110001111101110000 :
  (x[23:13] == 1989) ? 26'b10001001101111101111111100 :
  (x[23:13] == 1990) ? 26'b10001001101101100010001100 :
  (x[23:13] == 1991) ? 26'b10001001101011010100100000 :
  (x[23:13] == 1992) ? 26'b10001001101001000111000000 :
  (x[23:13] == 1993) ? 26'b10001001100110111001101000 :
  (x[23:13] == 1994) ? 26'b10001001100100101100010000 :
  (x[23:13] == 1995) ? 26'b10001001100010011111000100 :
  (x[23:13] == 1996) ? 26'b10001001100000010010000000 :
  (x[23:13] == 1997) ? 26'b10001001011110000101000000 :
  (x[23:13] == 1998) ? 26'b10001001011011111000000100 :
  (x[23:13] == 1999) ? 26'b10001001011001101011010000 :
  (x[23:13] == 2000) ? 26'b10001001010111011110101000 :
  (x[23:13] == 2001) ? 26'b10001001010101010010000000 :
  (x[23:13] == 2002) ? 26'b10001001010011000101100100 :
  (x[23:13] == 2003) ? 26'b10001001010000111001001100 :
  (x[23:13] == 2004) ? 26'b10001001001110101100111100 :
  (x[23:13] == 2005) ? 26'b10001001001100100000110000 :
  (x[23:13] == 2006) ? 26'b10001001001010010100110000 :
  (x[23:13] == 2007) ? 26'b10001001001000001000110100 :
  (x[23:13] == 2008) ? 26'b10001001000101111100111100 :
  (x[23:13] == 2009) ? 26'b10001001000011110001001100 :
  (x[23:13] == 2010) ? 26'b10001001000001100101100100 :
  (x[23:13] == 2011) ? 26'b10001000111111011010000100 :
  (x[23:13] == 2012) ? 26'b10001000111101001110101000 :
  (x[23:13] == 2013) ? 26'b10001000111011000011010000 :
  (x[23:13] == 2014) ? 26'b10001000111000111000000100 :
  (x[23:13] == 2015) ? 26'b10001000110110101101000000 :
  (x[23:13] == 2016) ? 26'b10001000110100100001111100 :
  (x[23:13] == 2017) ? 26'b10001000110010010111000100 :
  (x[23:13] == 2018) ? 26'b10001000110000001100010000 :
  (x[23:13] == 2019) ? 26'b10001000101110000001100100 :
  (x[23:13] == 2020) ? 26'b10001000101011110110111100 :
  (x[23:13] == 2021) ? 26'b10001000101001101100011100 :
  (x[23:13] == 2022) ? 26'b10001000100111100010000100 :
  (x[23:13] == 2023) ? 26'b10001000100101010111110000 :
  (x[23:13] == 2024) ? 26'b10001000100011001101101000 :
  (x[23:13] == 2025) ? 26'b10001000100001000011100000 :
  (x[23:13] == 2026) ? 26'b10001000011110111001100000 :
  (x[23:13] == 2027) ? 26'b10001000011100101111101000 :
  (x[23:13] == 2028) ? 26'b10001000011010100101111000 :
  (x[23:13] == 2029) ? 26'b10001000011000011100001100 :
  (x[23:13] == 2030) ? 26'b10001000010110010010101000 :
  (x[23:13] == 2031) ? 26'b10001000010100001001001000 :
  (x[23:13] == 2032) ? 26'b10001000010001111111110000 :
  (x[23:13] == 2033) ? 26'b10001000001111110110100000 :
  (x[23:13] == 2034) ? 26'b10001000001101101101011000 :
  (x[23:13] == 2035) ? 26'b10001000001011100100010000 :
  (x[23:13] == 2036) ? 26'b10001000001001011011010100 :
  (x[23:13] == 2037) ? 26'b10001000000111010010011100 :
  (x[23:13] == 2038) ? 26'b10001000000101001001101000 :
  (x[23:13] == 2039) ? 26'b10001000000011000001000000 :
  (x[23:13] == 2040) ? 26'b10001000000000111000011100 :
  (x[23:13] == 2041) ? 26'b10000111111110110000000000 :
  (x[23:13] == 2042) ? 26'b10000111111100100111101000 :
  (x[23:13] == 2043) ? 26'b10000111111010011111011000 :
  (x[23:13] == 2044) ? 26'b10000111111000010111001100 :
  (x[23:13] == 2045) ? 26'b10000111110110001111001000 :
  (x[23:13] == 2046) ? 26'b10000111110100000111001000 :
  26'b10000111110001111111010100 ;
  


  
  assign cube =
  (x[23:13] == 0) ? 26'b01011010011100011000010000 :
  (x[23:13] == 1) ? 26'b01011010010011111010100000 :
  (x[23:13] == 2) ? 26'b01011010001011011110000100 :
  (x[23:13] == 3) ? 26'b01011010000011000011000000 :
  (x[23:13] == 4) ? 26'b01011001111010101001001110 :
  (x[23:13] == 5) ? 26'b01011001110010010000110000 :
  (x[23:13] == 6) ? 26'b01011001101001111001011110 :
  (x[23:13] == 7) ? 26'b01011001100001100011101010 :
  (x[23:13] == 8) ? 26'b01011001011001001111000000 :
  (x[23:13] == 9) ? 26'b01011001010000111011101110 :
  (x[23:13] == 10) ? 26'b01011001001000101001101100 :
  (x[23:13] == 11) ? 26'b01011001000000011000111110 :
  (x[23:13] == 12) ? 26'b01011000111000001001100010 :
  (x[23:13] == 13) ? 26'b01011000101111111011010110 :
  (x[23:13] == 14) ? 26'b01011000100111101110011000 :
  (x[23:13] == 15) ? 26'b01011000011111100010101100 :
  (x[23:13] == 16) ? 26'b01011000010111011000010100 :
  (x[23:13] == 17) ? 26'b01011000001111001111000110 :
  (x[23:13] == 18) ? 26'b01011000000111000111001100 :
  (x[23:13] == 19) ? 26'b01010111111111000000100010 :
  (x[23:13] == 20) ? 26'b01010111110110111011000110 :
  (x[23:13] == 21) ? 26'b01010111101110110110111010 :
  (x[23:13] == 22) ? 26'b01010111100110110100000010 :
  (x[23:13] == 23) ? 26'b01010111011110110010010100 :
  (x[23:13] == 24) ? 26'b01010111010110110001110010 :
  (x[23:13] == 25) ? 26'b01010111001110110010100000 :
  (x[23:13] == 26) ? 26'b01010111000110110100011010 :
  (x[23:13] == 27) ? 26'b01010110111110110111101000 :
  (x[23:13] == 28) ? 26'b01010110110110111011111110 :
  (x[23:13] == 29) ? 26'b01010110101111000001100010 :
  (x[23:13] == 30) ? 26'b01010110100111001000010100 :
  (x[23:13] == 31) ? 26'b01010110011111010000001100 :
  (x[23:13] == 32) ? 26'b01010110010111011001011000 :
  (x[23:13] == 33) ? 26'b01010110001111100011110000 :
  (x[23:13] == 34) ? 26'b01010110000111101111010000 :
  (x[23:13] == 35) ? 26'b01010101111111111011111100 :
  (x[23:13] == 36) ? 26'b01010101111000001001110110 :
  (x[23:13] == 37) ? 26'b01010101110000011000111010 :
  (x[23:13] == 38) ? 26'b01010101101000101001000110 :
  (x[23:13] == 39) ? 26'b01010101100000111010011110 :
  (x[23:13] == 40) ? 26'b01010101011001001101000000 :
  (x[23:13] == 41) ? 26'b01010101010001100000110000 :
  (x[23:13] == 42) ? 26'b01010101001001110101100110 :
  (x[23:13] == 43) ? 26'b01010101000010001011100110 :
  (x[23:13] == 44) ? 26'b01010100111010100010110010 :
  (x[23:13] == 45) ? 26'b01010100110010111011000100 :
  (x[23:13] == 46) ? 26'b01010100101011010100100010 :
  (x[23:13] == 47) ? 26'b01010100100011101111001010 :
  (x[23:13] == 48) ? 26'b01010100011100001010110110 :
  (x[23:13] == 49) ? 26'b01010100010100100111101000 :
  (x[23:13] == 50) ? 26'b01010100001101000101100100 :
  (x[23:13] == 51) ? 26'b01010100000101100100101100 :
  (x[23:13] == 52) ? 26'b01010011111110000100110110 :
  (x[23:13] == 53) ? 26'b01010011110110100110001100 :
  (x[23:13] == 54) ? 26'b01010011101111001000100110 :
  (x[23:13] == 55) ? 26'b01010011100111101100001010 :
  (x[23:13] == 56) ? 26'b01010011100000010000110010 :
  (x[23:13] == 57) ? 26'b01010011011000110110011110 :
  (x[23:13] == 58) ? 26'b01010011010001011101010100 :
  (x[23:13] == 59) ? 26'b01010011001010000101001100 :
  (x[23:13] == 60) ? 26'b01010011000010101110001110 :
  (x[23:13] == 61) ? 26'b01010010111011011000010100 :
  (x[23:13] == 62) ? 26'b01010010110100000011011100 :
  (x[23:13] == 63) ? 26'b01010010101100101111101110 :
  (x[23:13] == 64) ? 26'b01010010100101011101000010 :
  (x[23:13] == 65) ? 26'b01010010011110001011011010 :
  (x[23:13] == 66) ? 26'b01010010010110111010110110 :
  (x[23:13] == 67) ? 26'b01010010001111101011011000 :
  (x[23:13] == 68) ? 26'b01010010001000011100111100 :
  (x[23:13] == 69) ? 26'b01010010000001001111100100 :
  (x[23:13] == 70) ? 26'b01010001111010000011001110 :
  (x[23:13] == 71) ? 26'b01010001110010111000000000 :
  (x[23:13] == 72) ? 26'b01010001101011101101110100 :
  (x[23:13] == 73) ? 26'b01010001100100100100100100 :
  (x[23:13] == 74) ? 26'b01010001011101011100011100 :
  (x[23:13] == 75) ? 26'b01010001010110010101011010 :
  (x[23:13] == 76) ? 26'b01010001001111001111010110 :
  (x[23:13] == 77) ? 26'b01010001001000001010010010 :
  (x[23:13] == 78) ? 26'b01010001000001000110010000 :
  (x[23:13] == 79) ? 26'b01010000111010000011010100 :
  (x[23:13] == 80) ? 26'b01010000110011000001010100 :
  (x[23:13] == 81) ? 26'b01010000101100000000011010 :
  (x[23:13] == 82) ? 26'b01010000100101000000011100 :
  (x[23:13] == 83) ? 26'b01010000011110000001100100 :
  (x[23:13] == 84) ? 26'b01010000010111000011101000 :
  (x[23:13] == 85) ? 26'b01010000010000000110110000 :
  (x[23:13] == 86) ? 26'b01010000001001001010110110 :
  (x[23:13] == 87) ? 26'b01010000000010001111111010 :
  (x[23:13] == 88) ? 26'b01001111111011010110000100 :
  (x[23:13] == 89) ? 26'b01001111110100011101001000 :
  (x[23:13] == 90) ? 26'b01001111101101100101001110 :
  (x[23:13] == 91) ? 26'b01001111100110101110010000 :
  (x[23:13] == 92) ? 26'b01001111011111111000010000 :
  (x[23:13] == 93) ? 26'b01001111011001000011010100 :
  (x[23:13] == 94) ? 26'b01001111010010001111010010 :
  (x[23:13] == 95) ? 26'b01001111001011011100001110 :
  (x[23:13] == 96) ? 26'b01001111000100101010001100 :
  (x[23:13] == 97) ? 26'b01001110111101111001000110 :
  (x[23:13] == 98) ? 26'b01001110110111001000111100 :
  (x[23:13] == 99) ? 26'b01001110110000011001110100 :
  (x[23:13] == 100) ? 26'b01001110101001101011101000 :
  (x[23:13] == 101) ? 26'b01001110100010111110010100 :
  (x[23:13] == 102) ? 26'b01001110011100010010000100 :
  (x[23:13] == 103) ? 26'b01001110010101100110101100 :
  (x[23:13] == 104) ? 26'b01001110001110111100001110 :
  (x[23:13] == 105) ? 26'b01001110001000010010110110 :
  (x[23:13] == 106) ? 26'b01001110000001101010010010 :
  (x[23:13] == 107) ? 26'b01001101111011000010110000 :
  (x[23:13] == 108) ? 26'b01001101110100011100000100 :
  (x[23:13] == 109) ? 26'b01001101101101110110011000 :
  (x[23:13] == 110) ? 26'b01001101100111010001100010 :
  (x[23:13] == 111) ? 26'b01001101100000101101101010 :
  (x[23:13] == 112) ? 26'b01001101011010001010110010 :
  (x[23:13] == 113) ? 26'b01001101010011101000110000 :
  (x[23:13] == 114) ? 26'b01001101001101000111100110 :
  (x[23:13] == 115) ? 26'b01001101000110100111011010 :
  (x[23:13] == 116) ? 26'b01001101000000001000001010 :
  (x[23:13] == 117) ? 26'b01001100111001101001110010 :
  (x[23:13] == 118) ? 26'b01001100110011001100011000 :
  (x[23:13] == 119) ? 26'b01001100101100101111110100 :
  (x[23:13] == 120) ? 26'b01001100100110010100001000 :
  (x[23:13] == 121) ? 26'b01001100011111111001011000 :
  (x[23:13] == 122) ? 26'b01001100011001011111100100 :
  (x[23:13] == 123) ? 26'b01001100010011000110100010 :
  (x[23:13] == 124) ? 26'b01001100001100101110011110 :
  (x[23:13] == 125) ? 26'b01001100000110010111010100 :
  (x[23:13] == 126) ? 26'b01001100000000000001000010 :
  (x[23:13] == 127) ? 26'b01001011111001101011100110 :
  (x[23:13] == 128) ? 26'b01001011110011010111000000 :
  (x[23:13] == 129) ? 26'b01001011101101000011010110 :
  (x[23:13] == 130) ? 26'b01001011100110110000100100 :
  (x[23:13] == 131) ? 26'b01001011100000011110100110 :
  (x[23:13] == 132) ? 26'b01001011011010001101100110 :
  (x[23:13] == 133) ? 26'b01001011010011111101011000 :
  (x[23:13] == 134) ? 26'b01001011001101101110000100 :
  (x[23:13] == 135) ? 26'b01001011000111011111101010 :
  (x[23:13] == 136) ? 26'b01001011000001010010000000 :
  (x[23:13] == 137) ? 26'b01001010111011000101010010 :
  (x[23:13] == 138) ? 26'b01001010110100111001011000 :
  (x[23:13] == 139) ? 26'b01001010101110101110010100 :
  (x[23:13] == 140) ? 26'b01001010101000100100001010 :
  (x[23:13] == 141) ? 26'b01001010100010011010110000 :
  (x[23:13] == 142) ? 26'b01001010011100010010010010 :
  (x[23:13] == 143) ? 26'b01001010010110001010101010 :
  (x[23:13] == 144) ? 26'b01001010010000000011101110 :
  (x[23:13] == 145) ? 26'b01001010001001111101110000 :
  (x[23:13] == 146) ? 26'b01001010000011111000100100 :
  (x[23:13] == 147) ? 26'b01001001111101110100010100 :
  (x[23:13] == 148) ? 26'b01001001110111110000110010 :
  (x[23:13] == 149) ? 26'b01001001110001101110000100 :
  (x[23:13] == 150) ? 26'b01001001101011101100001110 :
  (x[23:13] == 151) ? 26'b01001001100101101011001110 :
  (x[23:13] == 152) ? 26'b01001001011111101010111110 :
  (x[23:13] == 153) ? 26'b01001001011001101011100010 :
  (x[23:13] == 154) ? 26'b01001001010011101101000000 :
  (x[23:13] == 155) ? 26'b01001001001101101111001110 :
  (x[23:13] == 156) ? 26'b01001001000111110010001110 :
  (x[23:13] == 157) ? 26'b01001001000001110110000010 :
  (x[23:13] == 158) ? 26'b01001000111011111010110000 :
  (x[23:13] == 159) ? 26'b01001000110110000000001100 :
  (x[23:13] == 160) ? 26'b01001000110000000110010110 :
  (x[23:13] == 161) ? 26'b01001000101010001101011000 :
  (x[23:13] == 162) ? 26'b01001000100100010101010000 :
  (x[23:13] == 163) ? 26'b01001000011110011101111010 :
  (x[23:13] == 164) ? 26'b01001000011000100111010010 :
  (x[23:13] == 165) ? 26'b01001000010010110001011100 :
  (x[23:13] == 166) ? 26'b01001000001100111100100000 :
  (x[23:13] == 167) ? 26'b01001000000111001000010000 :
  (x[23:13] == 168) ? 26'b01001000000001010100110000 :
  (x[23:13] == 169) ? 26'b01000111111011100010000110 :
  (x[23:13] == 170) ? 26'b01000111110101110000001100 :
  (x[23:13] == 171) ? 26'b01000111101111111111000010 :
  (x[23:13] == 172) ? 26'b01000111101010001110101100 :
  (x[23:13] == 173) ? 26'b01000111100100011111001000 :
  (x[23:13] == 174) ? 26'b01000111011110110000010010 :
  (x[23:13] == 175) ? 26'b01000111011001000010001110 :
  (x[23:13] == 176) ? 26'b01000111010011010100111100 :
  (x[23:13] == 177) ? 26'b01000111001101101000011100 :
  (x[23:13] == 178) ? 26'b01000111000111111100101010 :
  (x[23:13] == 179) ? 26'b01000111000010010001101000 :
  (x[23:13] == 180) ? 26'b01000110111100100111010100 :
  (x[23:13] == 181) ? 26'b01000110110110111101111000 :
  (x[23:13] == 182) ? 26'b01000110110001010101000010 :
  (x[23:13] == 183) ? 26'b01000110101011101101000100 :
  (x[23:13] == 184) ? 26'b01000110100110000101110010 :
  (x[23:13] == 185) ? 26'b01000110100000011111010000 :
  (x[23:13] == 186) ? 26'b01000110011010111001011100 :
  (x[23:13] == 187) ? 26'b01000110010101010100011010 :
  (x[23:13] == 188) ? 26'b01000110001111110000000010 :
  (x[23:13] == 189) ? 26'b01000110001010001100011100 :
  (x[23:13] == 190) ? 26'b01000110000100101001101000 :
  (x[23:13] == 191) ? 26'b01000101111111000111100000 :
  (x[23:13] == 192) ? 26'b01000101111001100110001000 :
  (x[23:13] == 193) ? 26'b01000101110100000101011100 :
  (x[23:13] == 194) ? 26'b01000101101110100101100010 :
  (x[23:13] == 195) ? 26'b01000101101001000110010010 :
  (x[23:13] == 196) ? 26'b01000101100011100111101110 :
  (x[23:13] == 197) ? 26'b01000101011110001010000000 :
  (x[23:13] == 198) ? 26'b01000101011000101100111000 :
  (x[23:13] == 199) ? 26'b01000101010011010000100000 :
  (x[23:13] == 200) ? 26'b01000101001101110100111100 :
  (x[23:13] == 201) ? 26'b01000101001000011001111010 :
  (x[23:13] == 202) ? 26'b01000101000010111111101110 :
  (x[23:13] == 203) ? 26'b01000100111101100110001010 :
  (x[23:13] == 204) ? 26'b01000100111000001101011010 :
  (x[23:13] == 205) ? 26'b01000100110010110101001110 :
  (x[23:13] == 206) ? 26'b01000100101101011101110100 :
  (x[23:13] == 207) ? 26'b01000100101000000111000100 :
  (x[23:13] == 208) ? 26'b01000100100010110001000100 :
  (x[23:13] == 209) ? 26'b01000100011101011011110000 :
  (x[23:13] == 210) ? 26'b01000100011000000111000100 :
  (x[23:13] == 211) ? 26'b01000100010010110011000100 :
  (x[23:13] == 212) ? 26'b01000100001101011111110010 :
  (x[23:13] == 213) ? 26'b01000100001000001101001100 :
  (x[23:13] == 214) ? 26'b01000100000010111011010110 :
  (x[23:13] == 215) ? 26'b01000011111101101010001000 :
  (x[23:13] == 216) ? 26'b01000011111000011001100010 :
  (x[23:13] == 217) ? 26'b01000011110011001001101100 :
  (x[23:13] == 218) ? 26'b01000011101101111010011110 :
  (x[23:13] == 219) ? 26'b01000011101000101011111110 :
  (x[23:13] == 220) ? 26'b01000011100011011110001010 :
  (x[23:13] == 221) ? 26'b01000011011110010000111110 :
  (x[23:13] == 222) ? 26'b01000011011001000100011100 :
  (x[23:13] == 223) ? 26'b01000011010011111000101000 :
  (x[23:13] == 224) ? 26'b01000011001110101101011010 :
  (x[23:13] == 225) ? 26'b01000011001001100010111000 :
  (x[23:13] == 226) ? 26'b01000011000100011001000010 :
  (x[23:13] == 227) ? 26'b01000010111111001111111010 :
  (x[23:13] == 228) ? 26'b01000010111010000111010110 :
  (x[23:13] == 229) ? 26'b01000010110100111111011010 :
  (x[23:13] == 230) ? 26'b01000010101111111000001110 :
  (x[23:13] == 231) ? 26'b01000010101010110001101010 :
  (x[23:13] == 232) ? 26'b01000010100101101011101100 :
  (x[23:13] == 233) ? 26'b01000010100000100110011010 :
  (x[23:13] == 234) ? 26'b01000010011011100001110010 :
  (x[23:13] == 235) ? 26'b01000010010110011101110010 :
  (x[23:13] == 236) ? 26'b01000010010001011010011100 :
  (x[23:13] == 237) ? 26'b01000010001100010111101110 :
  (x[23:13] == 238) ? 26'b01000010000111010101101010 :
  (x[23:13] == 239) ? 26'b01000010000010010100010010 :
  (x[23:13] == 240) ? 26'b01000001111101010011011110 :
  (x[23:13] == 241) ? 26'b01000001111000010011010010 :
  (x[23:13] == 242) ? 26'b01000001110011010011110000 :
  (x[23:13] == 243) ? 26'b01000001101110010100110100 :
  (x[23:13] == 244) ? 26'b01000001101001010110101000 :
  (x[23:13] == 245) ? 26'b01000001100100011000111110 :
  (x[23:13] == 246) ? 26'b01000001011111011011111100 :
  (x[23:13] == 247) ? 26'b01000001011010011111100010 :
  (x[23:13] == 248) ? 26'b01000001010101100011110010 :
  (x[23:13] == 249) ? 26'b01000001010000101000101000 :
  (x[23:13] == 250) ? 26'b01000001001011101110000110 :
  (x[23:13] == 251) ? 26'b01000001000110110100001000 :
  (x[23:13] == 252) ? 26'b01000001000001111010110110 :
  (x[23:13] == 253) ? 26'b01000000111101000010000110 :
  (x[23:13] == 254) ? 26'b01000000111000001010000100 :
  (x[23:13] == 255) ? 26'b01000000110011010010100100 :
  (x[23:13] == 256) ? 26'b01000000101110011011101100 :
  (x[23:13] == 257) ? 26'b01000000101001100101011100 :
  (x[23:13] == 258) ? 26'b01000000100100101111110010 :
  (x[23:13] == 259) ? 26'b01000000011111111010110010 :
  (x[23:13] == 260) ? 26'b01000000011011000110010100 :
  (x[23:13] == 261) ? 26'b01000000010110010010100000 :
  (x[23:13] == 262) ? 26'b01000000010001011111010000 :
  (x[23:13] == 263) ? 26'b01000000001100101100100110 :
  (x[23:13] == 264) ? 26'b01000000000111111010011110 :
  (x[23:13] == 265) ? 26'b01000000000011001001000100 :
  (x[23:13] == 266) ? 26'b00111111111110011000001010 :
  (x[23:13] == 267) ? 26'b00111111111001100111110111 :
  (x[23:13] == 268) ? 26'b00111111110100111000001100 :
  (x[23:13] == 269) ? 26'b00111111110000001001000011 :
  (x[23:13] == 270) ? 26'b00111111101011011010100000 :
  (x[23:13] == 271) ? 26'b00111111100110101100100100 :
  (x[23:13] == 272) ? 26'b00111111100001111111001111 :
  (x[23:13] == 273) ? 26'b00111111011101010010011011 :
  (x[23:13] == 274) ? 26'b00111111011000100110001111 :
  (x[23:13] == 275) ? 26'b00111111010011111010100111 :
  (x[23:13] == 276) ? 26'b00111111001111001111100111 :
  (x[23:13] == 277) ? 26'b00111111001010100101001001 :
  (x[23:13] == 278) ? 26'b00111111000101111011001100 :
  (x[23:13] == 279) ? 26'b00111111000001010001111001 :
  (x[23:13] == 280) ? 26'b00111110111100101001001001 :
  (x[23:13] == 281) ? 26'b00111110111000000000111111 :
  (x[23:13] == 282) ? 26'b00111110110011011001010110 :
  (x[23:13] == 283) ? 26'b00111110101110110010010010 :
  (x[23:13] == 284) ? 26'b00111110101010001011110000 :
  (x[23:13] == 285) ? 26'b00111110100101100101110011 :
  (x[23:13] == 286) ? 26'b00111110100001000000011101 :
  (x[23:13] == 287) ? 26'b00111110011100011011101000 :
  (x[23:13] == 288) ? 26'b00111110010111110111011001 :
  (x[23:13] == 289) ? 26'b00111110010011010011101111 :
  (x[23:13] == 290) ? 26'b00111110001110110000100110 :
  (x[23:13] == 291) ? 26'b00111110001010001101111101 :
  (x[23:13] == 292) ? 26'b00111110000101101011111010 :
  (x[23:13] == 293) ? 26'b00111110000001001010011110 :
  (x[23:13] == 294) ? 26'b00111101111100101001100000 :
  (x[23:13] == 295) ? 26'b00111101111000001001000101 :
  (x[23:13] == 296) ? 26'b00111101110011101001010010 :
  (x[23:13] == 297) ? 26'b00111101101111001001111100 :
  (x[23:13] == 298) ? 26'b00111101101010101011001100 :
  (x[23:13] == 299) ? 26'b00111101100110001101000000 :
  (x[23:13] == 300) ? 26'b00111101100001101111010100 :
  (x[23:13] == 301) ? 26'b00111101011101010010001001 :
  (x[23:13] == 302) ? 26'b00111101011000110101100010 :
  (x[23:13] == 303) ? 26'b00111101010100011001100001 :
  (x[23:13] == 304) ? 26'b00111101001111111101111011 :
  (x[23:13] == 305) ? 26'b00111101001011100010111111 :
  (x[23:13] == 306) ? 26'b00111101000111001000011111 :
  (x[23:13] == 307) ? 26'b00111101000010101110100010 :
  (x[23:13] == 308) ? 26'b00111100111110010101001010 :
  (x[23:13] == 309) ? 26'b00111100111001111100010011 :
  (x[23:13] == 310) ? 26'b00111100110101100011111010 :
  (x[23:13] == 311) ? 26'b00111100110001001100001000 :
  (x[23:13] == 312) ? 26'b00111100101100110100110100 :
  (x[23:13] == 313) ? 26'b00111100101000011110000000 :
  (x[23:13] == 314) ? 26'b00111100100100000111110000 :
  (x[23:13] == 315) ? 26'b00111100011111110010000001 :
  (x[23:13] == 316) ? 26'b00111100011011011100110000 :
  (x[23:13] == 317) ? 26'b00111100010111001000000101 :
  (x[23:13] == 318) ? 26'b00111100010010110011110111 :
  (x[23:13] == 319) ? 26'b00111100001110100000001010 :
  (x[23:13] == 320) ? 26'b00111100001010001101000001 :
  (x[23:13] == 321) ? 26'b00111100000101111010011000 :
  (x[23:13] == 322) ? 26'b00111100000001101000001110 :
  (x[23:13] == 323) ? 26'b00111011111101010110100110 :
  (x[23:13] == 324) ? 26'b00111011111001000101011011 :
  (x[23:13] == 325) ? 26'b00111011110100110100110010 :
  (x[23:13] == 326) ? 26'b00111011110000100100101110 :
  (x[23:13] == 327) ? 26'b00111011101100010101000100 :
  (x[23:13] == 328) ? 26'b00111011101000000101111101 :
  (x[23:13] == 329) ? 26'b00111011100011110111010110 :
  (x[23:13] == 330) ? 26'b00111011011111101001001110 :
  (x[23:13] == 331) ? 26'b00111011011011011011101000 :
  (x[23:13] == 332) ? 26'b00111011010111001110011110 :
  (x[23:13] == 333) ? 26'b00111011010011000001110110 :
  (x[23:13] == 334) ? 26'b00111011001110110101101110 :
  (x[23:13] == 335) ? 26'b00111011001010101010001001 :
  (x[23:13] == 336) ? 26'b00111011000110011110111101 :
  (x[23:13] == 337) ? 26'b00111011000010010100010100 :
  (x[23:13] == 338) ? 26'b00111010111110001010000110 :
  (x[23:13] == 339) ? 26'b00111010111010000000011100 :
  (x[23:13] == 340) ? 26'b00111010110101110111001111 :
  (x[23:13] == 341) ? 26'b00111010110001101110100101 :
  (x[23:13] == 342) ? 26'b00111010101101100110010101 :
  (x[23:13] == 343) ? 26'b00111010101001011110100101 :
  (x[23:13] == 344) ? 26'b00111010100101010111010110 :
  (x[23:13] == 345) ? 26'b00111010100001010000100110 :
  (x[23:13] == 346) ? 26'b00111010011101001010001110 :
  (x[23:13] == 347) ? 26'b00111010011001000100011011 :
  (x[23:13] == 348) ? 26'b00111010010100111111000101 :
  (x[23:13] == 349) ? 26'b00111010010000111010001110 :
  (x[23:13] == 350) ? 26'b00111010001100110101111000 :
  (x[23:13] == 351) ? 26'b00111010001000110001111100 :
  (x[23:13] == 352) ? 26'b00111010000100101110011110 :
  (x[23:13] == 353) ? 26'b00111010000000101011011111 :
  (x[23:13] == 354) ? 26'b00111001111100101001000001 :
  (x[23:13] == 355) ? 26'b00111001111000100110111101 :
  (x[23:13] == 356) ? 26'b00111001110100100101010111 :
  (x[23:13] == 357) ? 26'b00111001110000100100010010 :
  (x[23:13] == 358) ? 26'b00111001101100100011100111 :
  (x[23:13] == 359) ? 26'b00111001101000100011011110 :
  (x[23:13] == 360) ? 26'b00111001100100100011101110 :
  (x[23:13] == 361) ? 26'b00111001100000100100100000 :
  (x[23:13] == 362) ? 26'b00111001011100100101101100 :
  (x[23:13] == 363) ? 26'b00111001011000100111010101 :
  (x[23:13] == 364) ? 26'b00111001010100101001100000 :
  (x[23:13] == 365) ? 26'b00111001010000101100000011 :
  (x[23:13] == 366) ? 26'b00111001001100101111000100 :
  (x[23:13] == 367) ? 26'b00111001001000110010100111 :
  (x[23:13] == 368) ? 26'b00111001000100110110100011 :
  (x[23:13] == 369) ? 26'b00111001000000111010111011 :
  (x[23:13] == 370) ? 26'b00111000111100111111110001 :
  (x[23:13] == 371) ? 26'b00111000111001000101000100 :
  (x[23:13] == 372) ? 26'b00111000110101001010110101 :
  (x[23:13] == 373) ? 26'b00111000110001010001000010 :
  (x[23:13] == 374) ? 26'b00111000101101010111100111 :
  (x[23:13] == 375) ? 26'b00111000101001011110110000 :
  (x[23:13] == 376) ? 26'b00111000100101100110001111 :
  (x[23:13] == 377) ? 26'b00111000100001101110010000 :
  (x[23:13] == 378) ? 26'b00111000011101110110101001 :
  (x[23:13] == 379) ? 26'b00111000011001111111100001 :
  (x[23:13] == 380) ? 26'b00111000010110001000110011 :
  (x[23:13] == 381) ? 26'b00111000010010010010100011 :
  (x[23:13] == 382) ? 26'b00111000001110011100101100 :
  (x[23:13] == 383) ? 26'b00111000001010100111010101 :
  (x[23:13] == 384) ? 26'b00111000000110110010010110 :
  (x[23:13] == 385) ? 26'b00111000000010111101110100 :
  (x[23:13] == 386) ? 26'b00110111111111001001101111 :
  (x[23:13] == 387) ? 26'b00110111111011010110000101 :
  (x[23:13] == 388) ? 26'b00110111110111100010110100 :
  (x[23:13] == 389) ? 26'b00110111110011110000000101 :
  (x[23:13] == 390) ? 26'b00110111101111111101101100 :
  (x[23:13] == 391) ? 26'b00110111101100001011110001 :
  (x[23:13] == 392) ? 26'b00110111101000011010010001 :
  (x[23:13] == 393) ? 26'b00110111100100101001001010 :
  (x[23:13] == 394) ? 26'b00110111100000111000011110 :
  (x[23:13] == 395) ? 26'b00110111011101001000001111 :
  (x[23:13] == 396) ? 26'b00110111011001011000011100 :
  (x[23:13] == 397) ? 26'b00110111010101101001000001 :
  (x[23:13] == 398) ? 26'b00110111010001111010000110 :
  (x[23:13] == 399) ? 26'b00110111001110001011100011 :
  (x[23:13] == 400) ? 26'b00110111001010011101010111 :
  (x[23:13] == 401) ? 26'b00110111000110101111101100 :
  (x[23:13] == 402) ? 26'b00110111000011000010011001 :
  (x[23:13] == 403) ? 26'b00110110111111010101100000 :
  (x[23:13] == 404) ? 26'b00110110111011101001000000 :
  (x[23:13] == 405) ? 26'b00110110110111111100111100 :
  (x[23:13] == 406) ? 26'b00110110110100010001010100 :
  (x[23:13] == 407) ? 26'b00110110110000100110000110 :
  (x[23:13] == 408) ? 26'b00110110101100111011010001 :
  (x[23:13] == 409) ? 26'b00110110101001010000110111 :
  (x[23:13] == 410) ? 26'b00110110100101100110111000 :
  (x[23:13] == 411) ? 26'b00110110100001111101010001 :
  (x[23:13] == 412) ? 26'b00110110011110010100000110 :
  (x[23:13] == 413) ? 26'b00110110011010101011010001 :
  (x[23:13] == 414) ? 26'b00110110010111000010111001 :
  (x[23:13] == 415) ? 26'b00110110010011011010111011 :
  (x[23:13] == 416) ? 26'b00110110001111110011010101 :
  (x[23:13] == 417) ? 26'b00110110001100001100001001 :
  (x[23:13] == 418) ? 26'b00110110001000100101011010 :
  (x[23:13] == 419) ? 26'b00110110000100111111000001 :
  (x[23:13] == 420) ? 26'b00110110000001011001000011 :
  (x[23:13] == 421) ? 26'b00110101111101110011011100 :
  (x[23:13] == 422) ? 26'b00110101111010001110010010 :
  (x[23:13] == 423) ? 26'b00110101110110101001100001 :
  (x[23:13] == 424) ? 26'b00110101110011000101001000 :
  (x[23:13] == 425) ? 26'b00110101101111100001001001 :
  (x[23:13] == 426) ? 26'b00110101101011111101100001 :
  (x[23:13] == 427) ? 26'b00110101101000011010010101 :
  (x[23:13] == 428) ? 26'b00110101100100110111011111 :
  (x[23:13] == 429) ? 26'b00110101100001010101000100 :
  (x[23:13] == 430) ? 26'b00110101011101110011000100 :
  (x[23:13] == 431) ? 26'b00110101011010010001011010 :
  (x[23:13] == 432) ? 26'b00110101010110110000000111 :
  (x[23:13] == 433) ? 26'b00110101010011001111001111 :
  (x[23:13] == 434) ? 26'b00110101001111101110110001 :
  (x[23:13] == 435) ? 26'b00110101001100001110101011 :
  (x[23:13] == 436) ? 26'b00110101001000101110111010 :
  (x[23:13] == 437) ? 26'b00110101000101001111100100 :
  (x[23:13] == 438) ? 26'b00110101000001110000101001 :
  (x[23:13] == 439) ? 26'b00110100111110010010000011 :
  (x[23:13] == 440) ? 26'b00110100111010110011110101 :
  (x[23:13] == 441) ? 26'b00110100110111010110000000 :
  (x[23:13] == 442) ? 26'b00110100110011111000100010 :
  (x[23:13] == 443) ? 26'b00110100110000011011011111 :
  (x[23:13] == 444) ? 26'b00110100101100111110110110 :
  (x[23:13] == 445) ? 26'b00110100101001100010011111 :
  (x[23:13] == 446) ? 26'b00110100100110000110100010 :
  (x[23:13] == 447) ? 26'b00110100100010101010111111 :
  (x[23:13] == 448) ? 26'b00110100011111001111110010 :
  (x[23:13] == 449) ? 26'b00110100011011110101000001 :
  (x[23:13] == 450) ? 26'b00110100011000011010011111 :
  (x[23:13] == 451) ? 26'b00110100010101000000011110 :
  (x[23:13] == 452) ? 26'b00110100010001100110101101 :
  (x[23:13] == 453) ? 26'b00110100001110001101011011 :
  (x[23:13] == 454) ? 26'b00110100001010110100011010 :
  (x[23:13] == 455) ? 26'b00110100000111011011110101 :
  (x[23:13] == 456) ? 26'b00110100000100000011100100 :
  (x[23:13] == 457) ? 26'b00110100000000101011101101 :
  (x[23:13] == 458) ? 26'b00110011111101010100001100 :
  (x[23:13] == 459) ? 26'b00110011111001111101000001 :
  (x[23:13] == 460) ? 26'b00110011110110100110001111 :
  (x[23:13] == 461) ? 26'b00110011110011001111110100 :
  (x[23:13] == 462) ? 26'b00110011101111111001101111 :
  (x[23:13] == 463) ? 26'b00110011101100100100000010 :
  (x[23:13] == 464) ? 26'b00110011101001001110101011 :
  (x[23:13] == 465) ? 26'b00110011100101111001101110 :
  (x[23:13] == 466) ? 26'b00110011100010100101000011 :
  (x[23:13] == 467) ? 26'b00110011011111010000110101 :
  (x[23:13] == 468) ? 26'b00110011011011111100111000 :
  (x[23:13] == 469) ? 26'b00110011011000101001010101 :
  (x[23:13] == 470) ? 26'b00110011010101010110000111 :
  (x[23:13] == 471) ? 26'b00110011010010000011001110 :
  (x[23:13] == 472) ? 26'b00110011001110110000110000 :
  (x[23:13] == 473) ? 26'b00110011001011011110100011 :
  (x[23:13] == 474) ? 26'b00110011001000001100110011 :
  (x[23:13] == 475) ? 26'b00110011000100111011010011 :
  (x[23:13] == 476) ? 26'b00110011000001101010001110 :
  (x[23:13] == 477) ? 26'b00110010111110011001011101 :
  (x[23:13] == 478) ? 26'b00110010111011001001000010 :
  (x[23:13] == 479) ? 26'b00110010110111111000111100 :
  (x[23:13] == 480) ? 26'b00110010110100101001001111 :
  (x[23:13] == 481) ? 26'b00110010110001011001110111 :
  (x[23:13] == 482) ? 26'b00110010101110001010110101 :
  (x[23:13] == 483) ? 26'b00110010101010111100001010 :
  (x[23:13] == 484) ? 26'b00110010100111101101110010 :
  (x[23:13] == 485) ? 26'b00110010100100011111110011 :
  (x[23:13] == 486) ? 26'b00110010100001010010001000 :
  (x[23:13] == 487) ? 26'b00110010011110000100110101 :
  (x[23:13] == 488) ? 26'b00110010011010110111110100 :
  (x[23:13] == 489) ? 26'b00110010010111101011001100 :
  (x[23:13] == 490) ? 26'b00110010010100011110111010 :
  (x[23:13] == 491) ? 26'b00110010010001010010111010 :
  (x[23:13] == 492) ? 26'b00110010001110000111010001 :
  (x[23:13] == 493) ? 26'b00110010001010111100000000 :
  (x[23:13] == 494) ? 26'b00110010000111110000111111 :
  (x[23:13] == 495) ? 26'b00110010000100100110011000 :
  (x[23:13] == 496) ? 26'b00110010000001011100000101 :
  (x[23:13] == 497) ? 26'b00110001111110010010000111 :
  (x[23:13] == 498) ? 26'b00110001111011001000100010 :
  (x[23:13] == 499) ? 26'b00110001110111111111001100 :
  (x[23:13] == 500) ? 26'b00110001110100110110010000 :
  (x[23:13] == 501) ? 26'b00110001110001101101100101 :
  (x[23:13] == 502) ? 26'b00110001101110100101010000 :
  (x[23:13] == 503) ? 26'b00110001101011011101010010 :
  (x[23:13] == 504) ? 26'b00110001101000010101100111 :
  (x[23:13] == 505) ? 26'b00110001100101001110010101 :
  (x[23:13] == 506) ? 26'b00110001100010000111010011 :
  (x[23:13] == 507) ? 26'b00110001011111000000100110 :
  (x[23:13] == 508) ? 26'b00110001011011111010010000 :
  (x[23:13] == 509) ? 26'b00110001011000110100010000 :
  (x[23:13] == 510) ? 26'b00110001010101101110011111 :
  (x[23:13] == 511) ? 26'b00110001010010101001000111 :
  (x[23:13] == 512) ? 26'b00110001001111100100000011 :
  (x[23:13] == 513) ? 26'b00110001001100011111010100 :
  (x[23:13] == 514) ? 26'b00110001001001011010111000 :
  (x[23:13] == 515) ? 26'b00110001000110010110110000 :
  (x[23:13] == 516) ? 26'b00110001000011010010111101 :
  (x[23:13] == 517) ? 26'b00110001000000001111100010 :
  (x[23:13] == 518) ? 26'b00110000111101001100010110 :
  (x[23:13] == 519) ? 26'b00110000111010001001011111 :
  (x[23:13] == 520) ? 26'b00110000110111000111000000 :
  (x[23:13] == 521) ? 26'b00110000110100000100110001 :
  (x[23:13] == 522) ? 26'b00110000110001000010110101 :
  (x[23:13] == 523) ? 26'b00110000101110000001010011 :
  (x[23:13] == 524) ? 26'b00110000101010111111111111 :
  (x[23:13] == 525) ? 26'b00110000100111111111000011 :
  (x[23:13] == 526) ? 26'b00110000100100111110010111 :
  (x[23:13] == 527) ? 26'b00110000100001111110000100 :
  (x[23:13] == 528) ? 26'b00110000011110111110000000 :
  (x[23:13] == 529) ? 26'b00110000011011111110010100 :
  (x[23:13] == 530) ? 26'b00110000011000111110111000 :
  (x[23:13] == 531) ? 26'b00110000010101111111110011 :
  (x[23:13] == 532) ? 26'b00110000010011000000111110 :
  (x[23:13] == 533) ? 26'b00110000010000000010100001 :
  (x[23:13] == 534) ? 26'b00110000001101000100010011 :
  (x[23:13] == 535) ? 26'b00110000001010000110011101 :
  (x[23:13] == 536) ? 26'b00110000000111001000110111 :
  (x[23:13] == 537) ? 26'b00110000000100001011101000 :
  (x[23:13] == 538) ? 26'b00110000000001001110101001 :
  (x[23:13] == 539) ? 26'b00101111111110010001111101 :
  (x[23:13] == 540) ? 26'b00101111111011010101100100 :
  (x[23:13] == 541) ? 26'b00101111111000011001011111 :
  (x[23:13] == 542) ? 26'b00101111110101011101101111 :
  (x[23:13] == 543) ? 26'b00101111110010100010010000 :
  (x[23:13] == 544) ? 26'b00101111101111100111000110 :
  (x[23:13] == 545) ? 26'b00101111101100101100001111 :
  (x[23:13] == 546) ? 26'b00101111101001110001101011 :
  (x[23:13] == 547) ? 26'b00101111100110110111011011 :
  (x[23:13] == 548) ? 26'b00101111100011111101011001 :
  (x[23:13] == 549) ? 26'b00101111100001000011110000 :
  (x[23:13] == 550) ? 26'b00101111011110001010010110 :
  (x[23:13] == 551) ? 26'b00101111011011010001001111 :
  (x[23:13] == 552) ? 26'b00101111011000011000011111 :
  (x[23:13] == 553) ? 26'b00101111010101011111111110 :
  (x[23:13] == 554) ? 26'b00101111010010100111110000 :
  (x[23:13] == 555) ? 26'b00101111001111101111110010 :
  (x[23:13] == 556) ? 26'b00101111001100111000001010 :
  (x[23:13] == 557) ? 26'b00101111001010000000110110 :
  (x[23:13] == 558) ? 26'b00101111000111001001110001 :
  (x[23:13] == 559) ? 26'b00101111000100010010111111 :
  (x[23:13] == 560) ? 26'b00101111000001011100100100 :
  (x[23:13] == 561) ? 26'b00101110111110100110010100 :
  (x[23:13] == 562) ? 26'b00101110111011110000011010 :
  (x[23:13] == 563) ? 26'b00101110111000111010110101 :
  (x[23:13] == 564) ? 26'b00101110110110000101011101 :
  (x[23:13] == 565) ? 26'b00101110110011010000011101 :
  (x[23:13] == 566) ? 26'b00101110110000011011101100 :
  (x[23:13] == 567) ? 26'b00101110101101100111001110 :
  (x[23:13] == 568) ? 26'b00101110101010110011000010 :
  (x[23:13] == 569) ? 26'b00101110100111111111000101 :
  (x[23:13] == 570) ? 26'b00101110100101001011011111 :
  (x[23:13] == 571) ? 26'b00101110100010011000001000 :
  (x[23:13] == 572) ? 26'b00101110011111100101000100 :
  (x[23:13] == 573) ? 26'b00101110011100110010010010 :
  (x[23:13] == 574) ? 26'b00101110011001111111101111 :
  (x[23:13] == 575) ? 26'b00101110010111001101100011 :
  (x[23:13] == 576) ? 26'b00101110010100011011100110 :
  (x[23:13] == 577) ? 26'b00101110010001101001111011 :
  (x[23:13] == 578) ? 26'b00101110001110111000100011 :
  (x[23:13] == 579) ? 26'b00101110001100000111011001 :
  (x[23:13] == 580) ? 26'b00101110001001010110100011 :
  (x[23:13] == 581) ? 26'b00101110000110100101111110 :
  (x[23:13] == 582) ? 26'b00101110000011110101101100 :
  (x[23:13] == 583) ? 26'b00101110000001000101101101 :
  (x[23:13] == 584) ? 26'b00101101111110010101111100 :
  (x[23:13] == 585) ? 26'b00101101111011100110011110 :
  (x[23:13] == 586) ? 26'b00101101111000110111010010 :
  (x[23:13] == 587) ? 26'b00101101110110001000010101 :
  (x[23:13] == 588) ? 26'b00101101110011011001101101 :
  (x[23:13] == 589) ? 26'b00101101110000101011010101 :
  (x[23:13] == 590) ? 26'b00101101101101111101001100 :
  (x[23:13] == 591) ? 26'b00101101101011001111010111 :
  (x[23:13] == 592) ? 26'b00101101101000100001110010 :
  (x[23:13] == 593) ? 26'b00101101100101110100011111 :
  (x[23:13] == 594) ? 26'b00101101100011000111011011 :
  (x[23:13] == 595) ? 26'b00101101100000011010101000 :
  (x[23:13] == 596) ? 26'b00101101011101101110001000 :
  (x[23:13] == 597) ? 26'b00101101011011000001111001 :
  (x[23:13] == 598) ? 26'b00101101011000010101111010 :
  (x[23:13] == 599) ? 26'b00101101010101101010001101 :
  (x[23:13] == 600) ? 26'b00101101010010111110110000 :
  (x[23:13] == 601) ? 26'b00101101010000010011100100 :
  (x[23:13] == 602) ? 26'b00101101001101101000101001 :
  (x[23:13] == 603) ? 26'b00101101001010111101111111 :
  (x[23:13] == 604) ? 26'b00101101001000010011100101 :
  (x[23:13] == 605) ? 26'b00101101000101101001011100 :
  (x[23:13] == 606) ? 26'b00101101000010111111100110 :
  (x[23:13] == 607) ? 26'b00101101000000010101111101 :
  (x[23:13] == 608) ? 26'b00101100111101101100100111 :
  (x[23:13] == 609) ? 26'b00101100111011000011100010 :
  (x[23:13] == 610) ? 26'b00101100111000011010101011 :
  (x[23:13] == 611) ? 26'b00101100110101110010000111 :
  (x[23:13] == 612) ? 26'b00101100110011001001110100 :
  (x[23:13] == 613) ? 26'b00101100110000100001101111 :
  (x[23:13] == 614) ? 26'b00101100101101111001111100 :
  (x[23:13] == 615) ? 26'b00101100101011010010011000 :
  (x[23:13] == 616) ? 26'b00101100101000101011000100 :
  (x[23:13] == 617) ? 26'b00101100100110000100000011 :
  (x[23:13] == 618) ? 26'b00101100100011011101010000 :
  (x[23:13] == 619) ? 26'b00101100100000110110101110 :
  (x[23:13] == 620) ? 26'b00101100011110010000011010 :
  (x[23:13] == 621) ? 26'b00101100011011101010011000 :
  (x[23:13] == 622) ? 26'b00101100011001000100101000 :
  (x[23:13] == 623) ? 26'b00101100010110011111000101 :
  (x[23:13] == 624) ? 26'b00101100010011111001110101 :
  (x[23:13] == 625) ? 26'b00101100010001010100110010 :
  (x[23:13] == 626) ? 26'b00101100001110110000000001 :
  (x[23:13] == 627) ? 26'b00101100001100001011100001 :
  (x[23:13] == 628) ? 26'b00101100001001100111001111 :
  (x[23:13] == 629) ? 26'b00101100000111000011001110 :
  (x[23:13] == 630) ? 26'b00101100000100011111011100 :
  (x[23:13] == 631) ? 26'b00101100000001111011111010 :
  (x[23:13] == 632) ? 26'b00101011111111011000100111 :
  (x[23:13] == 633) ? 26'b00101011111100110101100101 :
  (x[23:13] == 634) ? 26'b00101011111010010010110000 :
  (x[23:13] == 635) ? 26'b00101011110111110000001101 :
  (x[23:13] == 636) ? 26'b00101011110101001101111100 :
  (x[23:13] == 637) ? 26'b00101011110010101011111001 :
  (x[23:13] == 638) ? 26'b00101011110000001010000010 :
  (x[23:13] == 639) ? 26'b00101011101101101000100001 :
  (x[23:13] == 640) ? 26'b00101011101011000111001001 :
  (x[23:13] == 641) ? 26'b00101011101000100110000011 :
  (x[23:13] == 642) ? 26'b00101011100110000101001111 :
  (x[23:13] == 643) ? 26'b00101011100011100100100111 :
  (x[23:13] == 644) ? 26'b00101011100001000100010001 :
  (x[23:13] == 645) ? 26'b00101011011110100100001001 :
  (x[23:13] == 646) ? 26'b00101011011100000100010001 :
  (x[23:13] == 647) ? 26'b00101011011001100100100111 :
  (x[23:13] == 648) ? 26'b00101011010111000101001111 :
  (x[23:13] == 649) ? 26'b00101011010100100110000011 :
  (x[23:13] == 650) ? 26'b00101011010010000111000101 :
  (x[23:13] == 651) ? 26'b00101011001111101000011001 :
  (x[23:13] == 652) ? 26'b00101011001101001001111100 :
  (x[23:13] == 653) ? 26'b00101011001010101011101101 :
  (x[23:13] == 654) ? 26'b00101011001000001101110001 :
  (x[23:13] == 655) ? 26'b00101011000101110000000001 :
  (x[23:13] == 656) ? 26'b00101011000011010010011110 :
  (x[23:13] == 657) ? 26'b00101011000000110101001100 :
  (x[23:13] == 658) ? 26'b00101010111110011000001011 :
  (x[23:13] == 659) ? 26'b00101010111011111011010100 :
  (x[23:13] == 660) ? 26'b00101010111001011110110001 :
  (x[23:13] == 661) ? 26'b00101010110111000010011001 :
  (x[23:13] == 662) ? 26'b00101010110100100110010100 :
  (x[23:13] == 663) ? 26'b00101010110010001010011001 :
  (x[23:13] == 664) ? 26'b00101010101111101110101110 :
  (x[23:13] == 665) ? 26'b00101010101101010011010101 :
  (x[23:13] == 666) ? 26'b00101010101010111000001001 :
  (x[23:13] == 667) ? 26'b00101010101000011101001001 :
  (x[23:13] == 668) ? 26'b00101010100110000010011100 :
  (x[23:13] == 669) ? 26'b00101010100011100111111011 :
  (x[23:13] == 670) ? 26'b00101010100001001101101010 :
  (x[23:13] == 671) ? 26'b00101010011110110011100110 :
  (x[23:13] == 672) ? 26'b00101010011100011001110000 :
  (x[23:13] == 673) ? 26'b00101010011010000000001010 :
  (x[23:13] == 674) ? 26'b00101010010111100110110001 :
  (x[23:13] == 675) ? 26'b00101010010101001101100110 :
  (x[23:13] == 676) ? 26'b00101010010010110100101011 :
  (x[23:13] == 677) ? 26'b00101010010000011100000001 :
  (x[23:13] == 678) ? 26'b00101010001110000011100100 :
  (x[23:13] == 679) ? 26'b00101010001011101011010011 :
  (x[23:13] == 680) ? 26'b00101010001001010011001111 :
  (x[23:13] == 681) ? 26'b00101010000110111011011100 :
  (x[23:13] == 682) ? 26'b00101010000100100011110110 :
  (x[23:13] == 683) ? 26'b00101010000010001100100000 :
  (x[23:13] == 684) ? 26'b00101001111111110101010111 :
  (x[23:13] == 685) ? 26'b00101001111101011110011011 :
  (x[23:13] == 686) ? 26'b00101001111011000111101111 :
  (x[23:13] == 687) ? 26'b00101001111000110001010001 :
  (x[23:13] == 688) ? 26'b00101001110110011010111111 :
  (x[23:13] == 689) ? 26'b00101001110100000100111101 :
  (x[23:13] == 690) ? 26'b00101001110001101111001000 :
  (x[23:13] == 691) ? 26'b00101001101111011001100100 :
  (x[23:13] == 692) ? 26'b00101001101101000100001101 :
  (x[23:13] == 693) ? 26'b00101001101010101111000010 :
  (x[23:13] == 694) ? 26'b00101001101000011010000011 :
  (x[23:13] == 695) ? 26'b00101001100110000101010101 :
  (x[23:13] == 696) ? 26'b00101001100011110000110100 :
  (x[23:13] == 697) ? 26'b00101001100001011100011111 :
  (x[23:13] == 698) ? 26'b00101001011111001000011010 :
  (x[23:13] == 699) ? 26'b00101001011100110100100011 :
  (x[23:13] == 700) ? 26'b00101001011010100000110111 :
  (x[23:13] == 701) ? 26'b00101001011000001101011101 :
  (x[23:13] == 702) ? 26'b00101001010101111010001110 :
  (x[23:13] == 703) ? 26'b00101001010011100111001100 :
  (x[23:13] == 704) ? 26'b00101001010001010100011011 :
  (x[23:13] == 705) ? 26'b00101001001111000001110101 :
  (x[23:13] == 706) ? 26'b00101001001100101111011101 :
  (x[23:13] == 707) ? 26'b00101001001010011101010000 :
  (x[23:13] == 708) ? 26'b00101001001000001011010100 :
  (x[23:13] == 709) ? 26'b00101001000101111001100101 :
  (x[23:13] == 710) ? 26'b00101001000011101000000001 :
  (x[23:13] == 711) ? 26'b00101001000001010110101010 :
  (x[23:13] == 712) ? 26'b00101000111111000101100100 :
  (x[23:13] == 713) ? 26'b00101000111100110100101001 :
  (x[23:13] == 714) ? 26'b00101000111010100011111111 :
  (x[23:13] == 715) ? 26'b00101000111000010011011110 :
  (x[23:13] == 716) ? 26'b00101000110110000011001100 :
  (x[23:13] == 717) ? 26'b00101000110011110011000111 :
  (x[23:13] == 718) ? 26'b00101000110001100011001110 :
  (x[23:13] == 719) ? 26'b00101000101111010011100101 :
  (x[23:13] == 720) ? 26'b00101000101101000100001000 :
  (x[23:13] == 721) ? 26'b00101000101010110100110111 :
  (x[23:13] == 722) ? 26'b00101000101000100101110011 :
  (x[23:13] == 723) ? 26'b00101000100110010110111110 :
  (x[23:13] == 724) ? 26'b00101000100100001000010011 :
  (x[23:13] == 725) ? 26'b00101000100001111001110111 :
  (x[23:13] == 726) ? 26'b00101000011111101011101011 :
  (x[23:13] == 727) ? 26'b00101000011101011101101000 :
  (x[23:13] == 728) ? 26'b00101000011011001111110011 :
  (x[23:13] == 729) ? 26'b00101000011001000010001100 :
  (x[23:13] == 730) ? 26'b00101000010110110100110001 :
  (x[23:13] == 731) ? 26'b00101000010100100111100001 :
  (x[23:13] == 732) ? 26'b00101000010010011010011111 :
  (x[23:13] == 733) ? 26'b00101000010000001101101011 :
  (x[23:13] == 734) ? 26'b00101000001110000001000100 :
  (x[23:13] == 735) ? 26'b00101000001011110100101000 :
  (x[23:13] == 736) ? 26'b00101000001001101000011001 :
  (x[23:13] == 737) ? 26'b00101000000111011100011010 :
  (x[23:13] == 738) ? 26'b00101000000101010000100011 :
  (x[23:13] == 739) ? 26'b00101000000011000100111100 :
  (x[23:13] == 740) ? 26'b00101000000000111001100000 :
  (x[23:13] == 741) ? 26'b00100111111110101110010000 :
  (x[23:13] == 742) ? 26'b00100111111100100011010000 :
  (x[23:13] == 743) ? 26'b00100111111010011000011001 :
  (x[23:13] == 744) ? 26'b00100111111000001101110001 :
  (x[23:13] == 745) ? 26'b00100111110110000011010110 :
  (x[23:13] == 746) ? 26'b00100111110011111001000101 :
  (x[23:13] == 747) ? 26'b00100111110001101111000001 :
  (x[23:13] == 748) ? 26'b00100111101111100101001001 :
  (x[23:13] == 749) ? 26'b00100111101101011011100000 :
  (x[23:13] == 750) ? 26'b00100111101011010010000011 :
  (x[23:13] == 751) ? 26'b00100111101001001000101110 :
  (x[23:13] == 752) ? 26'b00100111100110111111101001 :
  (x[23:13] == 753) ? 26'b00100111100100110110110000 :
  (x[23:13] == 754) ? 26'b00100111100010101110000110 :
  (x[23:13] == 755) ? 26'b00100111100000100101100100 :
  (x[23:13] == 756) ? 26'b00100111011110011101001111 :
  (x[23:13] == 757) ? 26'b00100111011100010101001000 :
  (x[23:13] == 758) ? 26'b00100111011010001101001101 :
  (x[23:13] == 759) ? 26'b00100111011000000101011110 :
  (x[23:13] == 760) ? 26'b00100111010101111101111010 :
  (x[23:13] == 761) ? 26'b00100111010011110110100011 :
  (x[23:13] == 762) ? 26'b00100111010001101111011000 :
  (x[23:13] == 763) ? 26'b00100111001111101000010111 :
  (x[23:13] == 764) ? 26'b00100111001101100001100111 :
  (x[23:13] == 765) ? 26'b00100111001011011010111110 :
  (x[23:13] == 766) ? 26'b00100111001001010100100100 :
  (x[23:13] == 767) ? 26'b00100111000111001110010110 :
  (x[23:13] == 768) ? 26'b00100111000101001000010001 :
  (x[23:13] == 769) ? 26'b00100111000011000010011010 :
  (x[23:13] == 770) ? 26'b00100111000000111100101111 :
  (x[23:13] == 771) ? 26'b00100110111110110111001111 :
  (x[23:13] == 772) ? 26'b00100110111100110001111110 :
  (x[23:13] == 773) ? 26'b00100110111010101100110111 :
  (x[23:13] == 774) ? 26'b00100110111000100111111010 :
  (x[23:13] == 775) ? 26'b00100110110110100011001101 :
  (x[23:13] == 776) ? 26'b00100110110100011110100110 :
  (x[23:13] == 777) ? 26'b00100110110010011010010000 :
  (x[23:13] == 778) ? 26'b00100110110000010110000010 :
  (x[23:13] == 779) ? 26'b00100110101110010010000001 :
  (x[23:13] == 780) ? 26'b00100110101100001110001110 :
  (x[23:13] == 781) ? 26'b00100110101010001010100010 :
  (x[23:13] == 782) ? 26'b00100110101000000111000100 :
  (x[23:13] == 783) ? 26'b00100110100110000011110011 :
  (x[23:13] == 784) ? 26'b00100110100100000000101101 :
  (x[23:13] == 785) ? 26'b00100110100001111101110010 :
  (x[23:13] == 786) ? 26'b00100110011111111011000011 :
  (x[23:13] == 787) ? 26'b00100110011101111000011111 :
  (x[23:13] == 788) ? 26'b00100110011011110110001010 :
  (x[23:13] == 789) ? 26'b00100110011001110011111101 :
  (x[23:13] == 790) ? 26'b00100110010111110001111010 :
  (x[23:13] == 791) ? 26'b00100110010101110000000100 :
  (x[23:13] == 792) ? 26'b00100110010011101110011001 :
  (x[23:13] == 793) ? 26'b00100110010001101100111100 :
  (x[23:13] == 794) ? 26'b00100110001111101011101000 :
  (x[23:13] == 795) ? 26'b00100110001101101010011111 :
  (x[23:13] == 796) ? 26'b00100110001011101001100100 :
  (x[23:13] == 797) ? 26'b00100110001001101000110001 :
  (x[23:13] == 798) ? 26'b00100110000111101000001010 :
  (x[23:13] == 799) ? 26'b00100110000101100111110001 :
  (x[23:13] == 800) ? 26'b00100110000011100111100000 :
  (x[23:13] == 801) ? 26'b00100110000001100111011111 :
  (x[23:13] == 802) ? 26'b00100101111111100111100100 :
  (x[23:13] == 803) ? 26'b00100101111101100111110101 :
  (x[23:13] == 804) ? 26'b00100101111011101000010101 :
  (x[23:13] == 805) ? 26'b00100101111001101000111011 :
  (x[23:13] == 806) ? 26'b00100101110111101001101110 :
  (x[23:13] == 807) ? 26'b00100101110101101010101111 :
  (x[23:13] == 808) ? 26'b00100101110011101011110111 :
  (x[23:13] == 809) ? 26'b00100101110001101101001011 :
  (x[23:13] == 810) ? 26'b00100101101111101110101101 :
  (x[23:13] == 811) ? 26'b00100101101101110000010111 :
  (x[23:13] == 812) ? 26'b00100101101011110010001100 :
  (x[23:13] == 813) ? 26'b00100101101001110100001101 :
  (x[23:13] == 814) ? 26'b00100101100111110110011000 :
  (x[23:13] == 815) ? 26'b00100101100101111000110010 :
  (x[23:13] == 816) ? 26'b00100101100011111011010100 :
  (x[23:13] == 817) ? 26'b00100101100001111110000000 :
  (x[23:13] == 818) ? 26'b00100101100000000000110111 :
  (x[23:13] == 819) ? 26'b00100101011110000011111001 :
  (x[23:13] == 820) ? 26'b00100101011100000111000111 :
  (x[23:13] == 821) ? 26'b00100101011010001010011100 :
  (x[23:13] == 822) ? 26'b00100101011000001101111111 :
  (x[23:13] == 823) ? 26'b00100101010110010001101110 :
  (x[23:13] == 824) ? 26'b00100101010100010101100111 :
  (x[23:13] == 825) ? 26'b00100101010010011001101000 :
  (x[23:13] == 826) ? 26'b00100101010000011101111000 :
  (x[23:13] == 827) ? 26'b00100101001110100010001110 :
  (x[23:13] == 828) ? 26'b00100101001100100110110100 :
  (x[23:13] == 829) ? 26'b00100101001010101011100000 :
  (x[23:13] == 830) ? 26'b00100101001000110000011011 :
  (x[23:13] == 831) ? 26'b00100101000110110101011101 :
  (x[23:13] == 832) ? 26'b00100101000100111010101010 :
  (x[23:13] == 833) ? 26'b00100101000011000000000010 :
  (x[23:13] == 834) ? 26'b00100101000001000101100101 :
  (x[23:13] == 835) ? 26'b00100100111111001011010011 :
  (x[23:13] == 836) ? 26'b00100100111101010001001001 :
  (x[23:13] == 837) ? 26'b00100100111011010111001100 :
  (x[23:13] == 838) ? 26'b00100100111001011101011010 :
  (x[23:13] == 839) ? 26'b00100100110111100011101111 :
  (x[23:13] == 840) ? 26'b00100100110101101010010011 :
  (x[23:13] == 841) ? 26'b00100100110011110000111110 :
  (x[23:13] == 842) ? 26'b00100100110001110111110100 :
  (x[23:13] == 843) ? 26'b00100100101111111110110101 :
  (x[23:13] == 844) ? 26'b00100100101110000110000001 :
  (x[23:13] == 845) ? 26'b00100100101100001101010111 :
  (x[23:13] == 846) ? 26'b00100100101010010100111000 :
  (x[23:13] == 847) ? 26'b00100100101000011100100000 :
  (x[23:13] == 848) ? 26'b00100100100110100100010101 :
  (x[23:13] == 849) ? 26'b00100100100100101100010011 :
  (x[23:13] == 850) ? 26'b00100100100010110100011011 :
  (x[23:13] == 851) ? 26'b00100100100000111100110001 :
  (x[23:13] == 852) ? 26'b00100100011111000101001111 :
  (x[23:13] == 853) ? 26'b00100100011101001101110100 :
  (x[23:13] == 854) ? 26'b00100100011011010110100110 :
  (x[23:13] == 855) ? 26'b00100100011001011111100100 :
  (x[23:13] == 856) ? 26'b00100100010111101000101000 :
  (x[23:13] == 857) ? 26'b00100100010101110001111000 :
  (x[23:13] == 858) ? 26'b00100100010011111011010100 :
  (x[23:13] == 859) ? 26'b00100100010010000100111001 :
  (x[23:13] == 860) ? 26'b00100100010000001110100100 :
  (x[23:13] == 861) ? 26'b00100100001110011000011110 :
  (x[23:13] == 862) ? 26'b00100100001100100010100010 :
  (x[23:13] == 863) ? 26'b00100100001010101100101101 :
  (x[23:13] == 864) ? 26'b00100100001000110111000011 :
  (x[23:13] == 865) ? 26'b00100100000111000001100011 :
  (x[23:13] == 866) ? 26'b00100100000101001100001101 :
  (x[23:13] == 867) ? 26'b00100100000011010111000011 :
  (x[23:13] == 868) ? 26'b00100100000001100001111111 :
  (x[23:13] == 869) ? 26'b00100011111111101101001001 :
  (x[23:13] == 870) ? 26'b00100011111101111000011011 :
  (x[23:13] == 871) ? 26'b00100011111100000011110110 :
  (x[23:13] == 872) ? 26'b00100011111010001111011101 :
  (x[23:13] == 873) ? 26'b00100011111000011011001100 :
  (x[23:13] == 874) ? 26'b00100011110110100111000100 :
  (x[23:13] == 875) ? 26'b00100011110100110011000111 :
  (x[23:13] == 876) ? 26'b00100011110010111111010110 :
  (x[23:13] == 877) ? 26'b00100011110001001011101010 :
  (x[23:13] == 878) ? 26'b00100011101111011000001010 :
  (x[23:13] == 879) ? 26'b00100011101101100100110110 :
  (x[23:13] == 880) ? 26'b00100011101011110001101001 :
  (x[23:13] == 881) ? 26'b00100011101001111110100101 :
  (x[23:13] == 882) ? 26'b00100011101000001011101101 :
  (x[23:13] == 883) ? 26'b00100011100110011000111110 :
  (x[23:13] == 884) ? 26'b00100011100100100110010111 :
  (x[23:13] == 885) ? 26'b00100011100010110011111101 :
  (x[23:13] == 886) ? 26'b00100011100001000001101010 :
  (x[23:13] == 887) ? 26'b00100011011111001111011110 :
  (x[23:13] == 888) ? 26'b00100011011101011101100000 :
  (x[23:13] == 889) ? 26'b00100011011011101011101100 :
  (x[23:13] == 890) ? 26'b00100011011001111001111110 :
  (x[23:13] == 891) ? 26'b00100011011000001000011100 :
  (x[23:13] == 892) ? 26'b00100011010110010111000010 :
  (x[23:13] == 893) ? 26'b00100011010100100101110000 :
  (x[23:13] == 894) ? 26'b00100011010010110100101010 :
  (x[23:13] == 895) ? 26'b00100011010001000011101100 :
  (x[23:13] == 896) ? 26'b00100011001111010010111001 :
  (x[23:13] == 897) ? 26'b00100011001101100010010000 :
  (x[23:13] == 898) ? 26'b00100011001011110001101110 :
  (x[23:13] == 899) ? 26'b00100011001010000001010110 :
  (x[23:13] == 900) ? 26'b00100011001000010001001000 :
  (x[23:13] == 901) ? 26'b00100011000110100001000100 :
  (x[23:13] == 902) ? 26'b00100011000100110001000111 :
  (x[23:13] == 903) ? 26'b00100011000011000001010101 :
  (x[23:13] == 904) ? 26'b00100011000001010001101100 :
  (x[23:13] == 905) ? 26'b00100010111111100010001101 :
  (x[23:13] == 906) ? 26'b00100010111101110010110110 :
  (x[23:13] == 907) ? 26'b00100010111100000011101000 :
  (x[23:13] == 908) ? 26'b00100010111010010100100100 :
  (x[23:13] == 909) ? 26'b00100010111000100101100111 :
  (x[23:13] == 910) ? 26'b00100010110110110110111000 :
  (x[23:13] == 911) ? 26'b00100010110101001000001111 :
  (x[23:13] == 912) ? 26'b00100010110011011001101101 :
  (x[23:13] == 913) ? 26'b00100010110001101011011010 :
  (x[23:13] == 914) ? 26'b00100010101111111101001011 :
  (x[23:13] == 915) ? 26'b00100010101110001111001000 :
  (x[23:13] == 916) ? 26'b00100010101100100001001110 :
  (x[23:13] == 917) ? 26'b00100010101010110011011010 :
  (x[23:13] == 918) ? 26'b00100010101001000101110010 :
  (x[23:13] == 919) ? 26'b00100010100111011000010001 :
  (x[23:13] == 920) ? 26'b00100010100101101010111001 :
  (x[23:13] == 921) ? 26'b00100010100011111101101011 :
  (x[23:13] == 922) ? 26'b00100010100010010000100110 :
  (x[23:13] == 923) ? 26'b00100010100000100011101011 :
  (x[23:13] == 924) ? 26'b00100010011110110110110111 :
  (x[23:13] == 925) ? 26'b00100010011101001010001110 :
  (x[23:13] == 926) ? 26'b00100010011011011101101101 :
  (x[23:13] == 927) ? 26'b00100010011001110001010011 :
  (x[23:13] == 928) ? 26'b00100010011000000101000011 :
  (x[23:13] == 929) ? 26'b00100010010110011000111101 :
  (x[23:13] == 930) ? 26'b00100010010100101101000010 :
  (x[23:13] == 931) ? 26'b00100010010011000001001100 :
  (x[23:13] == 932) ? 26'b00100010010001010101011110 :
  (x[23:13] == 933) ? 26'b00100010001111101001111100 :
  (x[23:13] == 934) ? 26'b00100010001101111110100000 :
  (x[23:13] == 935) ? 26'b00100010001100010011001111 :
  (x[23:13] == 936) ? 26'b00100010001010101000001000 :
  (x[23:13] == 937) ? 26'b00100010001000111101000111 :
  (x[23:13] == 938) ? 26'b00100010000111010010001111 :
  (x[23:13] == 939) ? 26'b00100010000101100111011111 :
  (x[23:13] == 940) ? 26'b00100010000011111100111000 :
  (x[23:13] == 941) ? 26'b00100010000010010010011011 :
  (x[23:13] == 942) ? 26'b00100010000000101000000111 :
  (x[23:13] == 943) ? 26'b00100001111110111101111011 :
  (x[23:13] == 944) ? 26'b00100001111101010011110111 :
  (x[23:13] == 945) ? 26'b00100001111011101001111011 :
  (x[23:13] == 946) ? 26'b00100001111010000000001011 :
  (x[23:13] == 947) ? 26'b00100001111000010110011111 :
  (x[23:13] == 948) ? 26'b00100001110110101100111111 :
  (x[23:13] == 949) ? 26'b00100001110101000011100110 :
  (x[23:13] == 950) ? 26'b00100001110011011010010111 :
  (x[23:13] == 951) ? 26'b00100001110001110001001110 :
  (x[23:13] == 952) ? 26'b00100001110000001000001111 :
  (x[23:13] == 953) ? 26'b00100001101110011111011001 :
  (x[23:13] == 954) ? 26'b00100001101100110110101010 :
  (x[23:13] == 955) ? 26'b00100001101011001110000101 :
  (x[23:13] == 956) ? 26'b00100001101001100101101000 :
  (x[23:13] == 957) ? 26'b00100001100111111101010011 :
  (x[23:13] == 958) ? 26'b00100001100110010101000111 :
  (x[23:13] == 959) ? 26'b00100001100100101101000010 :
  (x[23:13] == 960) ? 26'b00100001100011000101001010 :
  (x[23:13] == 961) ? 26'b00100001100001011101010100 :
  (x[23:13] == 962) ? 26'b00100001011111110101101011 :
  (x[23:13] == 963) ? 26'b00100001011110001110001000 :
  (x[23:13] == 964) ? 26'b00100001011100100110101101 :
  (x[23:13] == 965) ? 26'b00100001011010111111011010 :
  (x[23:13] == 966) ? 26'b00100001011001011000010001 :
  (x[23:13] == 967) ? 26'b00100001010111110001010001 :
  (x[23:13] == 968) ? 26'b00100001010110001010011001 :
  (x[23:13] == 969) ? 26'b00100001010100100011100110 :
  (x[23:13] == 970) ? 26'b00100001010010111101000000 :
  (x[23:13] == 971) ? 26'b00100001010001010110011101 :
  (x[23:13] == 972) ? 26'b00100001001111110000000111 :
  (x[23:13] == 973) ? 26'b00100001001110001001110111 :
  (x[23:13] == 974) ? 26'b00100001001100100011110000 :
  (x[23:13] == 975) ? 26'b00100001001010111101110000 :
  (x[23:13] == 976) ? 26'b00100001001001010111111010 :
  (x[23:13] == 977) ? 26'b00100001000111110010001001 :
  (x[23:13] == 978) ? 26'b00100001000110001100100010 :
  (x[23:13] == 979) ? 26'b00100001000100100111000100 :
  (x[23:13] == 980) ? 26'b00100001000011000001101101 :
  (x[23:13] == 981) ? 26'b00100001000001011100011111 :
  (x[23:13] == 982) ? 26'b00100000111111110111010111 :
  (x[23:13] == 983) ? 26'b00100000111110010010011001 :
  (x[23:13] == 984) ? 26'b00100000111100101101100000 :
  (x[23:13] == 985) ? 26'b00100000111011001000110010 :
  (x[23:13] == 986) ? 26'b00100000111001100100001100 :
  (x[23:13] == 987) ? 26'b00100000110111111111101101 :
  (x[23:13] == 988) ? 26'b00100000110110011011010111 :
  (x[23:13] == 989) ? 26'b00100000110100110111000111 :
  (x[23:13] == 990) ? 26'b00100000110011010011000001 :
  (x[23:13] == 991) ? 26'b00100000110001101111000100 :
  (x[23:13] == 992) ? 26'b00100000110000001011001110 :
  (x[23:13] == 993) ? 26'b00100000101110100111011101 :
  (x[23:13] == 994) ? 26'b00100000101101000011111001 :
  (x[23:13] == 995) ? 26'b00100000101011100000010111 :
  (x[23:13] == 996) ? 26'b00100000101001111101000010 :
  (x[23:13] == 997) ? 26'b00100000101000011001110000 :
  (x[23:13] == 998) ? 26'b00100000100110110110101011 :
  (x[23:13] == 999) ? 26'b00100000100101010011101100 :
  (x[23:13] == 1000) ? 26'b00100000100011110000110011 :
  (x[23:13] == 1001) ? 26'b00100000100010001110000010 :
  (x[23:13] == 1002) ? 26'b00100000100000101011011100 :
  (x[23:13] == 1003) ? 26'b00100000011111001000111011 :
  (x[23:13] == 1004) ? 26'b00100000011101100110100001 :
  (x[23:13] == 1005) ? 26'b00100000011100000100010010 :
  (x[23:13] == 1006) ? 26'b00100000011010100010000111 :
  (x[23:13] == 1007) ? 26'b00100000011001000000001000 :
  (x[23:13] == 1008) ? 26'b00100000010111011110001011 :
  (x[23:13] == 1009) ? 26'b00100000010101111100011100 :
  (x[23:13] == 1010) ? 26'b00100000010100011010101111 :
  (x[23:13] == 1011) ? 26'b00100000010010111001001111 :
  (x[23:13] == 1012) ? 26'b00100000010001010111110101 :
  (x[23:13] == 1013) ? 26'b00100000001111110110100000 :
  (x[23:13] == 1014) ? 26'b00100000001110010101010100 :
  (x[23:13] == 1015) ? 26'b00100000001100110100001111 :
  (x[23:13] == 1016) ? 26'b00100000001011010011010011 :
  (x[23:13] == 1017) ? 26'b00100000001001110010011111 :
  (x[23:13] == 1018) ? 26'b00100000001000010001110010 :
  (x[23:13] == 1019) ? 26'b00100000000110110001001011 :
  (x[23:13] == 1020) ? 26'b00100000000101010000101101 :
  (x[23:13] == 1021) ? 26'b00100000000011110000011000 :
  (x[23:13] == 1022) ? 26'b00100000000010010000001001 :
  (x[23:13] == 1023) ? 26'b00100000000000110000000000 :
  (x[23:13] == 1024) ? 26'b11111111110100000000011000 :
  (x[23:13] == 1025) ? 26'b11111111011100000100001000 :
  (x[23:13] == 1026) ? 26'b11111111000100001011101000 :
  (x[23:13] == 1027) ? 26'b11111110101100010110110100 :
  (x[23:13] == 1028) ? 26'b11111110010100100101110000 :
  (x[23:13] == 1029) ? 26'b11111101111100111000011100 :
  (x[23:13] == 1030) ? 26'b11111101100101001110100100 :
  (x[23:13] == 1031) ? 26'b11111101001101101000100000 :
  (x[23:13] == 1032) ? 26'b11111100110110000110010000 :
  (x[23:13] == 1033) ? 26'b11111100011110100111010100 :
  (x[23:13] == 1034) ? 26'b11111100000111001100010000 :
  (x[23:13] == 1035) ? 26'b11111011101111110100110000 :
  (x[23:13] == 1036) ? 26'b11111011011000100000111000 :
  (x[23:13] == 1037) ? 26'b11111011000001010000101000 :
  (x[23:13] == 1038) ? 26'b11111010101010000011110100 :
  (x[23:13] == 1039) ? 26'b11111010010010111010110000 :
  (x[23:13] == 1040) ? 26'b11111001111011110101000100 :
  (x[23:13] == 1041) ? 26'b11111001100100110011000000 :
  (x[23:13] == 1042) ? 26'b11111001001101110100100000 :
  (x[23:13] == 1043) ? 26'b11111000110110111001100000 :
  (x[23:13] == 1044) ? 26'b11111000100000000001111100 :
  (x[23:13] == 1045) ? 26'b11111000001001001110000000 :
  (x[23:13] == 1046) ? 26'b11110111110010011101100000 :
  (x[23:13] == 1047) ? 26'b11110111011011110000011000 :
  (x[23:13] == 1048) ? 26'b11110111000101000110110100 :
  (x[23:13] == 1049) ? 26'b11110110101110100000110000 :
  (x[23:13] == 1050) ? 26'b11110110010111111110001000 :
  (x[23:13] == 1051) ? 26'b11110110000001011110110100 :
  (x[23:13] == 1052) ? 26'b11110101101011000011000000 :
  (x[23:13] == 1053) ? 26'b11110101010100101010100100 :
  (x[23:13] == 1054) ? 26'b11110100111110010101100000 :
  (x[23:13] == 1055) ? 26'b11110100101000000011111100 :
  (x[23:13] == 1056) ? 26'b11110100010001110101100100 :
  (x[23:13] == 1057) ? 26'b11110011111011101010110000 :
  (x[23:13] == 1058) ? 26'b11110011100101100011010000 :
  (x[23:13] == 1059) ? 26'b11110011001111011110111000 :
  (x[23:13] == 1060) ? 26'b11110010111001011110000100 :
  (x[23:13] == 1061) ? 26'b11110010100011100000100000 :
  (x[23:13] == 1062) ? 26'b11110010001101100110010100 :
  (x[23:13] == 1063) ? 26'b11110001110111101111010000 :
  (x[23:13] == 1064) ? 26'b11110001100001111011101000 :
  (x[23:13] == 1065) ? 26'b11110001001100001011001000 :
  (x[23:13] == 1066) ? 26'b11110000110110011110001000 :
  (x[23:13] == 1067) ? 26'b11110000100000110100001000 :
  (x[23:13] == 1068) ? 26'b11110000001011001101100100 :
  (x[23:13] == 1069) ? 26'b11101111110101101010001000 :
  (x[23:13] == 1070) ? 26'b11101111100000001001111000 :
  (x[23:13] == 1071) ? 26'b11101111001010101100111100 :
  (x[23:13] == 1072) ? 26'b11101110110101010011001100 :
  (x[23:13] == 1073) ? 26'b11101110011111111100011100 :
  (x[23:13] == 1074) ? 26'b11101110001010101001001000 :
  (x[23:13] == 1075) ? 26'b11101101110101011000111100 :
  (x[23:13] == 1076) ? 26'b11101101100000001011101100 :
  (x[23:13] == 1077) ? 26'b11101101001011000001101100 :
  (x[23:13] == 1078) ? 26'b11101100110101111010111100 :
  (x[23:13] == 1079) ? 26'b11101100100000110111011000 :
  (x[23:13] == 1080) ? 26'b11101100001011110110101100 :
  (x[23:13] == 1081) ? 26'b11101011110110111001010100 :
  (x[23:13] == 1082) ? 26'b11101011100001111110110100 :
  (x[23:13] == 1083) ? 26'b11101011001101000111101100 :
  (x[23:13] == 1084) ? 26'b11101010111000010011011000 :
  (x[23:13] == 1085) ? 26'b11101010100011100010010000 :
  (x[23:13] == 1086) ? 26'b11101010001110110100010000 :
  (x[23:13] == 1087) ? 26'b11101001111010001001010100 :
  (x[23:13] == 1088) ? 26'b11101001100101100001010000 :
  (x[23:13] == 1089) ? 26'b11101001010000111100010000 :
  (x[23:13] == 1090) ? 26'b11101000111100011010011000 :
  (x[23:13] == 1091) ? 26'b11101000100111111011100000 :
  (x[23:13] == 1092) ? 26'b11101000010011011111100000 :
  (x[23:13] == 1093) ? 26'b11100111111111000110100000 :
  (x[23:13] == 1094) ? 26'b11100111101010110000101000 :
  (x[23:13] == 1095) ? 26'b11100111010110011101100100 :
  (x[23:13] == 1096) ? 26'b11100111000010001101100000 :
  (x[23:13] == 1097) ? 26'b11100110101110000000011100 :
  (x[23:13] == 1098) ? 26'b11100110011001110110010100 :
  (x[23:13] == 1099) ? 26'b11100110000101101111001000 :
  (x[23:13] == 1100) ? 26'b11100101110001101010110000 :
  (x[23:13] == 1101) ? 26'b11100101011101101001100100 :
  (x[23:13] == 1102) ? 26'b11100101001001101011000100 :
  (x[23:13] == 1103) ? 26'b11100100110101101111100000 :
  (x[23:13] == 1104) ? 26'b11100100100001110110110000 :
  (x[23:13] == 1105) ? 26'b11100100001110000001000000 :
  (x[23:13] == 1106) ? 26'b11100011111010001110000100 :
  (x[23:13] == 1107) ? 26'b11100011100110011110000100 :
  (x[23:13] == 1108) ? 26'b11100011010010110000101000 :
  (x[23:13] == 1109) ? 26'b11100010111111000110011000 :
  (x[23:13] == 1110) ? 26'b11100010101011011110110000 :
  (x[23:13] == 1111) ? 26'b11100010010111111010001100 :
  (x[23:13] == 1112) ? 26'b11100010000100011000001000 :
  (x[23:13] == 1113) ? 26'b11100001110000111001000100 :
  (x[23:13] == 1114) ? 26'b11100001011101011100111000 :
  (x[23:13] == 1115) ? 26'b11100001001010000011010100 :
  (x[23:13] == 1116) ? 26'b11100000110110101100101000 :
  (x[23:13] == 1117) ? 26'b11100000100011011000100100 :
  (x[23:13] == 1118) ? 26'b11100000010000000111010100 :
  (x[23:13] == 1119) ? 26'b11011111111100111000111000 :
  (x[23:13] == 1120) ? 26'b11011111101001101101001000 :
  (x[23:13] == 1121) ? 26'b11011111010110100100001100 :
  (x[23:13] == 1122) ? 26'b11011111000011011110000000 :
  (x[23:13] == 1123) ? 26'b11011110110000011010100000 :
  (x[23:13] == 1124) ? 26'b11011110011101011001100100 :
  (x[23:13] == 1125) ? 26'b11011110001010011011011100 :
  (x[23:13] == 1126) ? 26'b11011101110111100000001000 :
  (x[23:13] == 1127) ? 26'b11011101100100100111011000 :
  (x[23:13] == 1128) ? 26'b11011101010001110001010000 :
  (x[23:13] == 1129) ? 26'b11011100111110111101111000 :
  (x[23:13] == 1130) ? 26'b11011100101100001101000100 :
  (x[23:13] == 1131) ? 26'b11011100011001011111001000 :
  (x[23:13] == 1132) ? 26'b11011100000110110011101100 :
  (x[23:13] == 1133) ? 26'b11011011110100001010110100 :
  (x[23:13] == 1134) ? 26'b11011011100001100100110000 :
  (x[23:13] == 1135) ? 26'b11011011001111000001000100 :
  (x[23:13] == 1136) ? 26'b11011010111100100000001000 :
  (x[23:13] == 1137) ? 26'b11011010101010000001111000 :
  (x[23:13] == 1138) ? 26'b11011010010111100110000100 :
  (x[23:13] == 1139) ? 26'b11011010000101001100111100 :
  (x[23:13] == 1140) ? 26'b11011001110010110110010100 :
  (x[23:13] == 1141) ? 26'b11011001100000100010010100 :
  (x[23:13] == 1142) ? 26'b11011001001110010001000000 :
  (x[23:13] == 1143) ? 26'b11011000111100000010000100 :
  (x[23:13] == 1144) ? 26'b11011000101001110101110100 :
  (x[23:13] == 1145) ? 26'b11011000010111101011111100 :
  (x[23:13] == 1146) ? 26'b11011000000101100100101100 :
  (x[23:13] == 1147) ? 26'b11010111110011100000000000 :
  (x[23:13] == 1148) ? 26'b11010111100001011101101100 :
  (x[23:13] == 1149) ? 26'b11010111001111011110000000 :
  (x[23:13] == 1150) ? 26'b11010110111101100000110100 :
  (x[23:13] == 1151) ? 26'b11010110101011100110001100 :
  (x[23:13] == 1152) ? 26'b11010110011001101101110100 :
  (x[23:13] == 1153) ? 26'b11010110000111111000001100 :
  (x[23:13] == 1154) ? 26'b11010101110110000100111100 :
  (x[23:13] == 1155) ? 26'b11010101100100010100000100 :
  (x[23:13] == 1156) ? 26'b11010101010010100101110000 :
  (x[23:13] == 1157) ? 26'b11010101000000111001110100 :
  (x[23:13] == 1158) ? 26'b11010100101111010000010100 :
  (x[23:13] == 1159) ? 26'b11010100011101101001010100 :
  (x[23:13] == 1160) ? 26'b11010100001100000100111000 :
  (x[23:13] == 1161) ? 26'b11010011111010100010101000 :
  (x[23:13] == 1162) ? 26'b11010011101001000010110100 :
  (x[23:13] == 1163) ? 26'b11010011010111100101100000 :
  (x[23:13] == 1164) ? 26'b11010011000110001010011100 :
  (x[23:13] == 1165) ? 26'b11010010110100110010000000 :
  (x[23:13] == 1166) ? 26'b11010010100011011011110100 :
  (x[23:13] == 1167) ? 26'b11010010010010000111111100 :
  (x[23:13] == 1168) ? 26'b11010010000000110110101000 :
  (x[23:13] == 1169) ? 26'b11010001101111100111011000 :
  (x[23:13] == 1170) ? 26'b11010001011110011010110000 :
  (x[23:13] == 1171) ? 26'b11010001001101010000011000 :
  (x[23:13] == 1172) ? 26'b11010000111100001000011000 :
  (x[23:13] == 1173) ? 26'b11010000101011000010101100 :
  (x[23:13] == 1174) ? 26'b11010000011001111111010100 :
  (x[23:13] == 1175) ? 26'b11010000001000111110010000 :
  (x[23:13] == 1176) ? 26'b11001111110111111111100000 :
  (x[23:13] == 1177) ? 26'b11001111100111000011001000 :
  (x[23:13] == 1178) ? 26'b11001111010110001001000000 :
  (x[23:13] == 1179) ? 26'b11001111000101010001001000 :
  (x[23:13] == 1180) ? 26'b11001110110100011011100000 :
  (x[23:13] == 1181) ? 26'b11001110100011101000010000 :
  (x[23:13] == 1182) ? 26'b11001110010010110111010100 :
  (x[23:13] == 1183) ? 26'b11001110000010001000100000 :
  (x[23:13] == 1184) ? 26'b11001101110001011100001100 :
  (x[23:13] == 1185) ? 26'b11001101100000110001111000 :
  (x[23:13] == 1186) ? 26'b11001101010000001001111100 :
  (x[23:13] == 1187) ? 26'b11001100111111100100010000 :
  (x[23:13] == 1188) ? 26'b11001100101111000000101000 :
  (x[23:13] == 1189) ? 26'b11001100011110011111011100 :
  (x[23:13] == 1190) ? 26'b11001100001110000000011000 :
  (x[23:13] == 1191) ? 26'b11001011111101100011100000 :
  (x[23:13] == 1192) ? 26'b11001011101101001000111000 :
  (x[23:13] == 1193) ? 26'b11001011011100110000100100 :
  (x[23:13] == 1194) ? 26'b11001011001100011010001100 :
  (x[23:13] == 1195) ? 26'b11001010111100000110001000 :
  (x[23:13] == 1196) ? 26'b11001010101011110100010000 :
  (x[23:13] == 1197) ? 26'b11001010011011100100100000 :
  (x[23:13] == 1198) ? 26'b11001010001011010111001000 :
  (x[23:13] == 1199) ? 26'b11001001111011001011101100 :
  (x[23:13] == 1200) ? 26'b11001001101011000010101000 :
  (x[23:13] == 1201) ? 26'b11001001011010111011011100 :
  (x[23:13] == 1202) ? 26'b11001001001010110110100100 :
  (x[23:13] == 1203) ? 26'b11001000111010110011101100 :
  (x[23:13] == 1204) ? 26'b11001000101010110011001100 :
  (x[23:13] == 1205) ? 26'b11001000011010110100100100 :
  (x[23:13] == 1206) ? 26'b11001000001010111000001100 :
  (x[23:13] == 1207) ? 26'b11000111111010111101110100 :
  (x[23:13] == 1208) ? 26'b11000111101011000101101100 :
  (x[23:13] == 1209) ? 26'b11000111011011001111100100 :
  (x[23:13] == 1210) ? 26'b11000111001011011011101100 :
  (x[23:13] == 1211) ? 26'b11000110111011101001110000 :
  (x[23:13] == 1212) ? 26'b11000110101011111001111000 :
  (x[23:13] == 1213) ? 26'b11000110011100001100001000 :
  (x[23:13] == 1214) ? 26'b11000110001100100000100000 :
  (x[23:13] == 1215) ? 26'b11000101111100110110111000 :
  (x[23:13] == 1216) ? 26'b11000101101101001111010100 :
  (x[23:13] == 1217) ? 26'b11000101011101101001110000 :
  (x[23:13] == 1218) ? 26'b11000101001110000110010000 :
  (x[23:13] == 1219) ? 26'b11000100111110100100111000 :
  (x[23:13] == 1220) ? 26'b11000100101111000101100100 :
  (x[23:13] == 1221) ? 26'b11000100011111101000001000 :
  (x[23:13] == 1222) ? 26'b11000100010000001100110100 :
  (x[23:13] == 1223) ? 26'b11000100000000110011100100 :
  (x[23:13] == 1224) ? 26'b11000011110001011100001100 :
  (x[23:13] == 1225) ? 26'b11000011100010000110110100 :
  (x[23:13] == 1226) ? 26'b11000011010010110011100100 :
  (x[23:13] == 1227) ? 26'b11000011000011100010011000 :
  (x[23:13] == 1228) ? 26'b11000010110100010011000100 :
  (x[23:13] == 1229) ? 26'b11000010100101000101101000 :
  (x[23:13] == 1230) ? 26'b11000010010101111010011000 :
  (x[23:13] == 1231) ? 26'b11000010000110110000111000 :
  (x[23:13] == 1232) ? 26'b11000001110111101001100000 :
  (x[23:13] == 1233) ? 26'b11000001101000100100000100 :
  (x[23:13] == 1234) ? 26'b11000001011001100000100000 :
  (x[23:13] == 1235) ? 26'b11000001001010011110111100 :
  (x[23:13] == 1236) ? 26'b11000000111011011111011000 :
  (x[23:13] == 1237) ? 26'b11000000101100100001110000 :
  (x[23:13] == 1238) ? 26'b11000000011101100101111100 :
  (x[23:13] == 1239) ? 26'b11000000001110101100001000 :
  (x[23:13] == 1240) ? 26'b10111111111111110100011000 :
  (x[23:13] == 1241) ? 26'b10111111110000111110010000 :
  (x[23:13] == 1242) ? 26'b10111111100010001010010000 :
  (x[23:13] == 1243) ? 26'b10111111010011011000000100 :
  (x[23:13] == 1244) ? 26'b10111111000100100111110000 :
  (x[23:13] == 1245) ? 26'b10111110110101111001100000 :
  (x[23:13] == 1246) ? 26'b10111110100111001100111100 :
  (x[23:13] == 1247) ? 26'b10111110011000100010011000 :
  (x[23:13] == 1248) ? 26'b10111110001001111001101100 :
  (x[23:13] == 1249) ? 26'b10111101111011010010110000 :
  (x[23:13] == 1250) ? 26'b10111101101100101101110100 :
  (x[23:13] == 1251) ? 26'b10111101011110001010110100 :
  (x[23:13] == 1252) ? 26'b10111101001111101001100000 :
  (x[23:13] == 1253) ? 26'b10111101000001001010001000 :
  (x[23:13] == 1254) ? 26'b10111100110010101100101000 :
  (x[23:13] == 1255) ? 26'b10111100100100010000111000 :
  (x[23:13] == 1256) ? 26'b10111100010101110111000100 :
  (x[23:13] == 1257) ? 26'b10111100000111011110111100 :
  (x[23:13] == 1258) ? 26'b10111011111001001000110000 :
  (x[23:13] == 1259) ? 26'b10111011101010110100011000 :
  (x[23:13] == 1260) ? 26'b10111011011100100001110000 :
  (x[23:13] == 1261) ? 26'b10111011001110010001001000 :
  (x[23:13] == 1262) ? 26'b10111011000000000010001000 :
  (x[23:13] == 1263) ? 26'b10111010110001110101000100 :
  (x[23:13] == 1264) ? 26'b10111010100011101001101000 :
  (x[23:13] == 1265) ? 26'b10111010010101100000000100 :
  (x[23:13] == 1266) ? 26'b10111010000111011000011000 :
  (x[23:13] == 1267) ? 26'b10111001111001010010011000 :
  (x[23:13] == 1268) ? 26'b10111001101011001110001100 :
  (x[23:13] == 1269) ? 26'b10111001011101001011101000 :
  (x[23:13] == 1270) ? 26'b10111001001111001011000000 :
  (x[23:13] == 1271) ? 26'b10111001000001001100000100 :
  (x[23:13] == 1272) ? 26'b10111000110011001110111100 :
  (x[23:13] == 1273) ? 26'b10111000100101010011100100 :
  (x[23:13] == 1274) ? 26'b10111000010111011010000000 :
  (x[23:13] == 1275) ? 26'b10111000001001100010000100 :
  (x[23:13] == 1276) ? 26'b10110111111011101011110100 :
  (x[23:13] == 1277) ? 26'b10110111101101110111011100 :
  (x[23:13] == 1278) ? 26'b10110111100000000100101000 :
  (x[23:13] == 1279) ? 26'b10110111010010010011110000 :
  (x[23:13] == 1280) ? 26'b10110111000100100100100000 :
  (x[23:13] == 1281) ? 26'b10110110110110110110111000 :
  (x[23:13] == 1282) ? 26'b10110110101001001011000100 :
  (x[23:13] == 1283) ? 26'b10110110011011100000111100 :
  (x[23:13] == 1284) ? 26'b10110110001101111000101000 :
  (x[23:13] == 1285) ? 26'b10110110000000010001110000 :
  (x[23:13] == 1286) ? 26'b10110101110010101100111000 :
  (x[23:13] == 1287) ? 26'b10110101100101001001100100 :
  (x[23:13] == 1288) ? 26'b10110101010111100111101100 :
  (x[23:13] == 1289) ? 26'b10110101001010000111110100 :
  (x[23:13] == 1290) ? 26'b10110100111100101001011100 :
  (x[23:13] == 1291) ? 26'b10110100101111001100110100 :
  (x[23:13] == 1292) ? 26'b10110100100001110001110100 :
  (x[23:13] == 1293) ? 26'b10110100010100011000011100 :
  (x[23:13] == 1294) ? 26'b10110100000111000000111000 :
  (x[23:13] == 1295) ? 26'b10110011111001101010110000 :
  (x[23:13] == 1296) ? 26'b10110011101100010110100000 :
  (x[23:13] == 1297) ? 26'b10110011011111000011110000 :
  (x[23:13] == 1298) ? 26'b10110011010001110010101000 :
  (x[23:13] == 1299) ? 26'b10110011000100100011001000 :
  (x[23:13] == 1300) ? 26'b10110010110111010101010100 :
  (x[23:13] == 1301) ? 26'b10110010101010001001001000 :
  (x[23:13] == 1302) ? 26'b10110010011100111110100000 :
  (x[23:13] == 1303) ? 26'b10110010001111110101101000 :
  (x[23:13] == 1304) ? 26'b10110010000010101110001100 :
  (x[23:13] == 1305) ? 26'b10110001110101101000011100 :
  (x[23:13] == 1306) ? 26'b10110001101000100100011000 :
  (x[23:13] == 1307) ? 26'b10110001011011100001110100 :
  (x[23:13] == 1308) ? 26'b10110001001110100000110100 :
  (x[23:13] == 1309) ? 26'b10110001000001100001011100 :
  (x[23:13] == 1310) ? 26'b10110000110100100011110000 :
  (x[23:13] == 1311) ? 26'b10110000100111100111100000 :
  (x[23:13] == 1312) ? 26'b10110000011010101100111000 :
  (x[23:13] == 1313) ? 26'b10110000001101110011110100 :
  (x[23:13] == 1314) ? 26'b10110000000000111100010100 :
  (x[23:13] == 1315) ? 26'b10101111110100000110011100 :
  (x[23:13] == 1316) ? 26'b10101111100111010010000100 :
  (x[23:13] == 1317) ? 26'b10101111011010011111010100 :
  (x[23:13] == 1318) ? 26'b10101111001101101110000100 :
  (x[23:13] == 1319) ? 26'b10101111000000111110010100 :
  (x[23:13] == 1320) ? 26'b10101110110100010000010000 :
  (x[23:13] == 1321) ? 26'b10101110100111100011101000 :
  (x[23:13] == 1322) ? 26'b10101110011010111000011100 :
  (x[23:13] == 1323) ? 26'b10101110001110001110111100 :
  (x[23:13] == 1324) ? 26'b10101110000001100110111100 :
  (x[23:13] == 1325) ? 26'b10101101110101000000011100 :
  (x[23:13] == 1326) ? 26'b10101101101000011011011100 :
  (x[23:13] == 1327) ? 26'b10101101011011111000000000 :
  (x[23:13] == 1328) ? 26'b10101101001111010110000100 :
  (x[23:13] == 1329) ? 26'b10101101000010110101100100 :
  (x[23:13] == 1330) ? 26'b10101100110110010110101000 :
  (x[23:13] == 1331) ? 26'b10101100101001111001010000 :
  (x[23:13] == 1332) ? 26'b10101100011101011101010000 :
  (x[23:13] == 1333) ? 26'b10101100010001000010111000 :
  (x[23:13] == 1334) ? 26'b10101100000100101001110100 :
  (x[23:13] == 1335) ? 26'b10101011111000010010011100 :
  (x[23:13] == 1336) ? 26'b10101011101011111100011100 :
  (x[23:13] == 1337) ? 26'b10101011011111100111111000 :
  (x[23:13] == 1338) ? 26'b10101011010011010100110100 :
  (x[23:13] == 1339) ? 26'b10101011000111000011010100 :
  (x[23:13] == 1340) ? 26'b10101010111010110011000100 :
  (x[23:13] == 1341) ? 26'b10101010101110100100100100 :
  (x[23:13] == 1342) ? 26'b10101010100010010111011000 :
  (x[23:13] == 1343) ? 26'b10101010010110001011101000 :
  (x[23:13] == 1344) ? 26'b10101010001010000001001100 :
  (x[23:13] == 1345) ? 26'b10101001111101111000010100 :
  (x[23:13] == 1346) ? 26'b10101001110001110001000100 :
  (x[23:13] == 1347) ? 26'b10101001100101101011001000 :
  (x[23:13] == 1348) ? 26'b10101001011001100110100100 :
  (x[23:13] == 1349) ? 26'b10101001001101100011011000 :
  (x[23:13] == 1350) ? 26'b10101001000001100001101100 :
  (x[23:13] == 1351) ? 26'b10101000110101100001100100 :
  (x[23:13] == 1352) ? 26'b10101000101001100010101100 :
  (x[23:13] == 1353) ? 26'b10101000011101100101001100 :
  (x[23:13] == 1354) ? 26'b10101000010001101001001100 :
  (x[23:13] == 1355) ? 26'b10101000000101101110101000 :
  (x[23:13] == 1356) ? 26'b10100111111001110101011000 :
  (x[23:13] == 1357) ? 26'b10100111101101111101101100 :
  (x[23:13] == 1358) ? 26'b10100111100010000111011000 :
  (x[23:13] == 1359) ? 26'b10100111010110010010010000 :
  (x[23:13] == 1360) ? 26'b10100111001010011110101100 :
  (x[23:13] == 1361) ? 26'b10100110111110101100100000 :
  (x[23:13] == 1362) ? 26'b10100110110010111011101100 :
  (x[23:13] == 1363) ? 26'b10100110100111001100001100 :
  (x[23:13] == 1364) ? 26'b10100110011011011110000100 :
  (x[23:13] == 1365) ? 26'b10100110001111110001011100 :
  (x[23:13] == 1366) ? 26'b10100110000100000110001000 :
  (x[23:13] == 1367) ? 26'b10100101111000011100000100 :
  (x[23:13] == 1368) ? 26'b10100101101100110011011100 :
  (x[23:13] == 1369) ? 26'b10100101100001001100010000 :
  (x[23:13] == 1370) ? 26'b10100101010101100110011000 :
  (x[23:13] == 1371) ? 26'b10100101001010000001110100 :
  (x[23:13] == 1372) ? 26'b10100100111110011110101000 :
  (x[23:13] == 1373) ? 26'b10100100110010111100110100 :
  (x[23:13] == 1374) ? 26'b10100100100111011100010100 :
  (x[23:13] == 1375) ? 26'b10100100011011111101000100 :
  (x[23:13] == 1376) ? 26'b10100100010000011111010100 :
  (x[23:13] == 1377) ? 26'b10100100000101000010111000 :
  (x[23:13] == 1378) ? 26'b10100011111001100111101000 :
  (x[23:13] == 1379) ? 26'b10100011101110001101110100 :
  (x[23:13] == 1380) ? 26'b10100011100010110101010100 :
  (x[23:13] == 1381) ? 26'b10100011010111011110000000 :
  (x[23:13] == 1382) ? 26'b10100011001100001000001000 :
  (x[23:13] == 1383) ? 26'b10100011000000110011100100 :
  (x[23:13] == 1384) ? 26'b10100010110101100000010000 :
  (x[23:13] == 1385) ? 26'b10100010101010001110011100 :
  (x[23:13] == 1386) ? 26'b10100010011110111101101100 :
  (x[23:13] == 1387) ? 26'b10100010010011101110011000 :
  (x[23:13] == 1388) ? 26'b10100010001000100000001000 :
  (x[23:13] == 1389) ? 26'b10100001111101010011100000 :
  (x[23:13] == 1390) ? 26'b10100001110010001000000000 :
  (x[23:13] == 1391) ? 26'b10100001100110111101110000 :
  (x[23:13] == 1392) ? 26'b10100001011011110100110100 :
  (x[23:13] == 1393) ? 26'b10100001010000101101001100 :
  (x[23:13] == 1394) ? 26'b10100001000101100110110000 :
  (x[23:13] == 1395) ? 26'b10100000111010100001101100 :
  (x[23:13] == 1396) ? 26'b10100000101111011101111000 :
  (x[23:13] == 1397) ? 26'b10100000100100011011010100 :
  (x[23:13] == 1398) ? 26'b10100000011001011010001000 :
  (x[23:13] == 1399) ? 26'b10100000001110011010000100 :
  (x[23:13] == 1400) ? 26'b10100000000011011011001100 :
  (x[23:13] == 1401) ? 26'b10011111111000011101101100 :
  (x[23:13] == 1402) ? 26'b10011111101101100001100000 :
  (x[23:13] == 1403) ? 26'b10011111100010100110011100 :
  (x[23:13] == 1404) ? 26'b10011111010111101100100100 :
  (x[23:13] == 1405) ? 26'b10011111001100110100000100 :
  (x[23:13] == 1406) ? 26'b10011111000001111100101100 :
  (x[23:13] == 1407) ? 26'b10011110110111000110101000 :
  (x[23:13] == 1408) ? 26'b10011110101100010001110100 :
  (x[23:13] == 1409) ? 26'b10011110100001011110010000 :
  (x[23:13] == 1410) ? 26'b10011110010110101011111000 :
  (x[23:13] == 1411) ? 26'b10011110001011111010101000 :
  (x[23:13] == 1412) ? 26'b10011110000001001010110000 :
  (x[23:13] == 1413) ? 26'b10011101110110011100000000 :
  (x[23:13] == 1414) ? 26'b10011101101011101110011100 :
  (x[23:13] == 1415) ? 26'b10011101100001000010001000 :
  (x[23:13] == 1416) ? 26'b10011101010110010111000000 :
  (x[23:13] == 1417) ? 26'b10011101001011101101001100 :
  (x[23:13] == 1418) ? 26'b10011101000001000100100100 :
  (x[23:13] == 1419) ? 26'b10011100110110011101000100 :
  (x[23:13] == 1420) ? 26'b10011100101011110110101100 :
  (x[23:13] == 1421) ? 26'b10011100100001010001100100 :
  (x[23:13] == 1422) ? 26'b10011100010110101101101100 :
  (x[23:13] == 1423) ? 26'b10011100001100001010111000 :
  (x[23:13] == 1424) ? 26'b10011100000001101001011100 :
  (x[23:13] == 1425) ? 26'b10011011110111001000111100 :
  (x[23:13] == 1426) ? 26'b10011011101100101001111000 :
  (x[23:13] == 1427) ? 26'b10011011100010001011111000 :
  (x[23:13] == 1428) ? 26'b10011011010111101110111100 :
  (x[23:13] == 1429) ? 26'b10011011001101010011010100 :
  (x[23:13] == 1430) ? 26'b10011011000010111000110100 :
  (x[23:13] == 1431) ? 26'b10011010111000011111011100 :
  (x[23:13] == 1432) ? 26'b10011010101110000111011000 :
  (x[23:13] == 1433) ? 26'b10011010100011110000010100 :
  (x[23:13] == 1434) ? 26'b10011010011001011010100000 :
  (x[23:13] == 1435) ? 26'b10011010001111000101110000 :
  (x[23:13] == 1436) ? 26'b10011010000100110010001100 :
  (x[23:13] == 1437) ? 26'b10011001111010011111110000 :
  (x[23:13] == 1438) ? 26'b10011001110000001110011100 :
  (x[23:13] == 1439) ? 26'b10011001100101111110011000 :
  (x[23:13] == 1440) ? 26'b10011001011011101111010100 :
  (x[23:13] == 1441) ? 26'b10011001010001100001100000 :
  (x[23:13] == 1442) ? 26'b10011001000111010100110100 :
  (x[23:13] == 1443) ? 26'b10011000111101001001010000 :
  (x[23:13] == 1444) ? 26'b10011000110010111110110100 :
  (x[23:13] == 1445) ? 26'b10011000101000110101011100 :
  (x[23:13] == 1446) ? 26'b10011000011110101101001100 :
  (x[23:13] == 1447) ? 26'b10011000010100100110000100 :
  (x[23:13] == 1448) ? 26'b10011000001010100000000100 :
  (x[23:13] == 1449) ? 26'b10011000000000011011001100 :
  (x[23:13] == 1450) ? 26'b10010111110110010111100000 :
  (x[23:13] == 1451) ? 26'b10010111101100010100110100 :
  (x[23:13] == 1452) ? 26'b10010111100010010011001100 :
  (x[23:13] == 1453) ? 26'b10010111011000010010111000 :
  (x[23:13] == 1454) ? 26'b10010111001110010011100000 :
  (x[23:13] == 1455) ? 26'b10010111000100010101001100 :
  (x[23:13] == 1456) ? 26'b10010110111010011000001100 :
  (x[23:13] == 1457) ? 26'b10010110110000011100000100 :
  (x[23:13] == 1458) ? 26'b10010110100110100001000100 :
  (x[23:13] == 1459) ? 26'b10010110011100100111001100 :
  (x[23:13] == 1460) ? 26'b10010110010010101110100000 :
  (x[23:13] == 1461) ? 26'b10010110001000110110110000 :
  (x[23:13] == 1462) ? 26'b10010101111111000000001000 :
  (x[23:13] == 1463) ? 26'b10010101110101001010100100 :
  (x[23:13] == 1464) ? 26'b10010101101011010110001000 :
  (x[23:13] == 1465) ? 26'b10010101100001100010101000 :
  (x[23:13] == 1466) ? 26'b10010101010111110000010100 :
  (x[23:13] == 1467) ? 26'b10010101001101111111001000 :
  (x[23:13] == 1468) ? 26'b10010101000100001110110100 :
  (x[23:13] == 1469) ? 26'b10010100111010011111101100 :
  (x[23:13] == 1470) ? 26'b10010100110000110001101100 :
  (x[23:13] == 1471) ? 26'b10010100100111000100101100 :
  (x[23:13] == 1472) ? 26'b10010100011101011000110000 :
  (x[23:13] == 1473) ? 26'b10010100010011101101101100 :
  (x[23:13] == 1474) ? 26'b10010100001010000011111000 :
  (x[23:13] == 1475) ? 26'b10010100000000011011000000 :
  (x[23:13] == 1476) ? 26'b10010011110110110011010000 :
  (x[23:13] == 1477) ? 26'b10010011101101001100011100 :
  (x[23:13] == 1478) ? 26'b10010011100011100110110000 :
  (x[23:13] == 1479) ? 26'b10010011011010000010001100 :
  (x[23:13] == 1480) ? 26'b10010011010000011110100000 :
  (x[23:13] == 1481) ? 26'b10010011000110111011111000 :
  (x[23:13] == 1482) ? 26'b10010010111101011010010100 :
  (x[23:13] == 1483) ? 26'b10010010110011111001110100 :
  (x[23:13] == 1484) ? 26'b10010010101010011010010100 :
  (x[23:13] == 1485) ? 26'b10010010100000111011110000 :
  (x[23:13] == 1486) ? 26'b10010010010111011110010100 :
  (x[23:13] == 1487) ? 26'b10010010001110000001111000 :
  (x[23:13] == 1488) ? 26'b10010010000100100110011000 :
  (x[23:13] == 1489) ? 26'b10010001111011001011111100 :
  (x[23:13] == 1490) ? 26'b10010001110001110010100100 :
  (x[23:13] == 1491) ? 26'b10010001101000011010010000 :
  (x[23:13] == 1492) ? 26'b10010001011111000010111000 :
  (x[23:13] == 1493) ? 26'b10010001010101101100100000 :
  (x[23:13] == 1494) ? 26'b10010001001100010111000000 :
  (x[23:13] == 1495) ? 26'b10010001000011000010100100 :
  (x[23:13] == 1496) ? 26'b10010000111001101111001100 :
  (x[23:13] == 1497) ? 26'b10010000110000011100110000 :
  (x[23:13] == 1498) ? 26'b10010000100111001011011100 :
  (x[23:13] == 1499) ? 26'b10010000011101111010111100 :
  (x[23:13] == 1500) ? 26'b10010000010100101011100000 :
  (x[23:13] == 1501) ? 26'b10010000001011011101000100 :
  (x[23:13] == 1502) ? 26'b10010000000010001111100100 :
  (x[23:13] == 1503) ? 26'b10001111111001000011000100 :
  (x[23:13] == 1504) ? 26'b10001111101111110111100000 :
  (x[23:13] == 1505) ? 26'b10001111100110101100111100 :
  (x[23:13] == 1506) ? 26'b10001111011101100011011000 :
  (x[23:13] == 1507) ? 26'b10001111010100011010110100 :
  (x[23:13] == 1508) ? 26'b10001111001011010011001100 :
  (x[23:13] == 1509) ? 26'b10001111000010001100100100 :
  (x[23:13] == 1510) ? 26'b10001110111001000110111000 :
  (x[23:13] == 1511) ? 26'b10001110110000000010000000 :
  (x[23:13] == 1512) ? 26'b10001110100110111110011000 :
  (x[23:13] == 1513) ? 26'b10001110011101111011100100 :
  (x[23:13] == 1514) ? 26'b10001110010100111001101100 :
  (x[23:13] == 1515) ? 26'b10001110001011111000110000 :
  (x[23:13] == 1516) ? 26'b10001110000010111000110000 :
  (x[23:13] == 1517) ? 26'b10001101111001111001110000 :
  (x[23:13] == 1518) ? 26'b10001101110000111011101100 :
  (x[23:13] == 1519) ? 26'b10001101100111111110100100 :
  (x[23:13] == 1520) ? 26'b10001101011111000010011000 :
  (x[23:13] == 1521) ? 26'b10001101010110000111001100 :
  (x[23:13] == 1522) ? 26'b10001101001101001100110100 :
  (x[23:13] == 1523) ? 26'b10001101000100010011100000 :
  (x[23:13] == 1524) ? 26'b10001100111011011011000100 :
  (x[23:13] == 1525) ? 26'b10001100110010100011100000 :
  (x[23:13] == 1526) ? 26'b10001100101001101100111100 :
  (x[23:13] == 1527) ? 26'b10001100100000110111010100 :
  (x[23:13] == 1528) ? 26'b10001100011000000010101000 :
  (x[23:13] == 1529) ? 26'b10001100001111001110110000 :
  (x[23:13] == 1530) ? 26'b10001100000110011011111100 :
  (x[23:13] == 1531) ? 26'b10001011111101101010000000 :
  (x[23:13] == 1532) ? 26'b10001011110100111000111100 :
  (x[23:13] == 1533) ? 26'b10001011101100001000110100 :
  (x[23:13] == 1534) ? 26'b10001011100011011001100100 :
  (x[23:13] == 1535) ? 26'b10001011011010101011010100 :
  (x[23:13] == 1536) ? 26'b10001011010001111101110100 :
  (x[23:13] == 1537) ? 26'b10001011001001010001011100 :
  (x[23:13] == 1538) ? 26'b10001011000000100101110000 :
  (x[23:13] == 1539) ? 26'b10001010110111111011001000 :
  (x[23:13] == 1540) ? 26'b10001010101111010001010100 :
  (x[23:13] == 1541) ? 26'b10001010100110101000100000 :
  (x[23:13] == 1542) ? 26'b10001010011110000000100000 :
  (x[23:13] == 1543) ? 26'b10001010010101011001011100 :
  (x[23:13] == 1544) ? 26'b10001010001100110011001100 :
  (x[23:13] == 1545) ? 26'b10001010000100001101111000 :
  (x[23:13] == 1546) ? 26'b10001001111011101001011100 :
  (x[23:13] == 1547) ? 26'b10001001110011000101111000 :
  (x[23:13] == 1548) ? 26'b10001001101010100011010000 :
  (x[23:13] == 1549) ? 26'b10001001100010000001100000 :
  (x[23:13] == 1550) ? 26'b10001001011001100000100100 :
  (x[23:13] == 1551) ? 26'b10001001010001000000100000 :
  (x[23:13] == 1552) ? 26'b10001001001000100001011100 :
  (x[23:13] == 1553) ? 26'b10001001000000000011001100 :
  (x[23:13] == 1554) ? 26'b10001000110111100101110000 :
  (x[23:13] == 1555) ? 26'b10001000101111001001010000 :
  (x[23:13] == 1556) ? 26'b10001000100110101101101000 :
  (x[23:13] == 1557) ? 26'b10001000011110010010110000 :
  (x[23:13] == 1558) ? 26'b10001000010101111000110100 :
  (x[23:13] == 1559) ? 26'b10001000001101011111111000 :
  (x[23:13] == 1560) ? 26'b10001000000101000111101000 :
  (x[23:13] == 1561) ? 26'b10000111111100110000001100 :
  (x[23:13] == 1562) ? 26'b10000111110100011001110000 :
  (x[23:13] == 1563) ? 26'b10000111101100000100001000 :
  (x[23:13] == 1564) ? 26'b10000111100011101111010100 :
  (x[23:13] == 1565) ? 26'b10000111011011011011011000 :
  (x[23:13] == 1566) ? 26'b10000111010011001000011000 :
  (x[23:13] == 1567) ? 26'b10000111001010110110000100 :
  (x[23:13] == 1568) ? 26'b10000111000010100100110000 :
  (x[23:13] == 1569) ? 26'b10000110111010010100010000 :
  (x[23:13] == 1570) ? 26'b10000110110010000100011000 :
  (x[23:13] == 1571) ? 26'b10000110101001110101100000 :
  (x[23:13] == 1572) ? 26'b10000110100001100111101000 :
  (x[23:13] == 1573) ? 26'b10000110011001011010011000 :
  (x[23:13] == 1574) ? 26'b10000110010001001110000000 :
  (x[23:13] == 1575) ? 26'b10000110001001000010100000 :
  (x[23:13] == 1576) ? 26'b10000110000000110111110100 :
  (x[23:13] == 1577) ? 26'b10000101111000101101111100 :
  (x[23:13] == 1578) ? 26'b10000101110000100100110100 :
  (x[23:13] == 1579) ? 26'b10000101101000011100101000 :
  (x[23:13] == 1580) ? 26'b10000101100000010101010000 :
  (x[23:13] == 1581) ? 26'b10000101011000001110101100 :
  (x[23:13] == 1582) ? 26'b10000101010000001000111100 :
  (x[23:13] == 1583) ? 26'b10000101001000000100000000 :
  (x[23:13] == 1584) ? 26'b10000100111111111111111000 :
  (x[23:13] == 1585) ? 26'b10000100110111111100100100 :
  (x[23:13] == 1586) ? 26'b10000100101111111010001000 :
  (x[23:13] == 1587) ? 26'b10000100100111111000011000 :
  (x[23:13] == 1588) ? 26'b10000100011111110111100000 :
  (x[23:13] == 1589) ? 26'b10000100010111110111011100 :
  (x[23:13] == 1590) ? 26'b10000100001111111000001000 :
  (x[23:13] == 1591) ? 26'b10000100000111111001101100 :
  (x[23:13] == 1592) ? 26'b10000011111111111100000000 :
  (x[23:13] == 1593) ? 26'b10000011110111111111001100 :
  (x[23:13] == 1594) ? 26'b10000011110000000011000100 :
  (x[23:13] == 1595) ? 26'b10000011101000000111110100 :
  (x[23:13] == 1596) ? 26'b10000011100000001101011000 :
  (x[23:13] == 1597) ? 26'b10000011011000010011101100 :
  (x[23:13] == 1598) ? 26'b10000011010000011010110100 :
  (x[23:13] == 1599) ? 26'b10000011001000100010101000 :
  (x[23:13] == 1600) ? 26'b10000011000000101011011000 :
  (x[23:13] == 1601) ? 26'b10000010111000110100111000 :
  (x[23:13] == 1602) ? 26'b10000010110000111111000100 :
  (x[23:13] == 1603) ? 26'b10000010101001001010001000 :
  (x[23:13] == 1604) ? 26'b10000010100001010101111100 :
  (x[23:13] == 1605) ? 26'b10000010011001100010011100 :
  (x[23:13] == 1606) ? 26'b10000010010001101111111100 :
  (x[23:13] == 1607) ? 26'b10000010001001111110000100 :
  (x[23:13] == 1608) ? 26'b10000010000010001101000000 :
  (x[23:13] == 1609) ? 26'b10000001111010011100100100 :
  (x[23:13] == 1610) ? 26'b10000001110010101101000100 :
  (x[23:13] == 1611) ? 26'b10000001101010111110011000 :
  (x[23:13] == 1612) ? 26'b10000001100011010000010100 :
  (x[23:13] == 1613) ? 26'b10000001011011100011001100 :
  (x[23:13] == 1614) ? 26'b10000001010011110110101100 :
  (x[23:13] == 1615) ? 26'b10000001001100001010111100 :
  (x[23:13] == 1616) ? 26'b10000001000100011111111100 :
  (x[23:13] == 1617) ? 26'b10000000111100110101110000 :
  (x[23:13] == 1618) ? 26'b10000000110101001100011000 :
  (x[23:13] == 1619) ? 26'b10000000101101100011101100 :
  (x[23:13] == 1620) ? 26'b10000000100101111011101100 :
  (x[23:13] == 1621) ? 26'b10000000011110010100100100 :
  (x[23:13] == 1622) ? 26'b10000000010110101110001100 :
  (x[23:13] == 1623) ? 26'b10000000001111001000011100 :
  (x[23:13] == 1624) ? 26'b10000000000111100011101000 :
  (x[23:13] == 1625) ? 26'b01111111111111111111011010 :
  (x[23:13] == 1626) ? 26'b01111111111000011011111110 :
  (x[23:13] == 1627) ? 26'b01111111110000111001001110 :
  (x[23:13] == 1628) ? 26'b01111111101001010111010100 :
  (x[23:13] == 1629) ? 26'b01111111100001110110000100 :
  (x[23:13] == 1630) ? 26'b01111111011010010101100110 :
  (x[23:13] == 1631) ? 26'b01111111010010110101111000 :
  (x[23:13] == 1632) ? 26'b01111111001011010110110100 :
  (x[23:13] == 1633) ? 26'b01111111000011111000100100 :
  (x[23:13] == 1634) ? 26'b01111110111100011011000000 :
  (x[23:13] == 1635) ? 26'b01111110110100111110001110 :
  (x[23:13] == 1636) ? 26'b01111110101101100010001000 :
  (x[23:13] == 1637) ? 26'b01111110100110000110110000 :
  (x[23:13] == 1638) ? 26'b01111110011110101100001000 :
  (x[23:13] == 1639) ? 26'b01111110010111010010010000 :
  (x[23:13] == 1640) ? 26'b01111110001111111001000110 :
  (x[23:13] == 1641) ? 26'b01111110001000100000101000 :
  (x[23:13] == 1642) ? 26'b01111110000001001000110100 :
  (x[23:13] == 1643) ? 26'b01111101111001110001111000 :
  (x[23:13] == 1644) ? 26'b01111101110010011011100100 :
  (x[23:13] == 1645) ? 26'b01111101101011000101111000 :
  (x[23:13] == 1646) ? 26'b01111101100011110000111100 :
  (x[23:13] == 1647) ? 26'b01111101011100011100110010 :
  (x[23:13] == 1648) ? 26'b01111101010101001001011000 :
  (x[23:13] == 1649) ? 26'b01111101001101110110100110 :
  (x[23:13] == 1650) ? 26'b01111101000110100100100110 :
  (x[23:13] == 1651) ? 26'b01111100111111010011010010 :
  (x[23:13] == 1652) ? 26'b01111100111000000010100110 :
  (x[23:13] == 1653) ? 26'b01111100110000110010101100 :
  (x[23:13] == 1654) ? 26'b01111100101001100011011100 :
  (x[23:13] == 1655) ? 26'b01111100100010010100110110 :
  (x[23:13] == 1656) ? 26'b01111100011011000111000100 :
  (x[23:13] == 1657) ? 26'b01111100010011111001111010 :
  (x[23:13] == 1658) ? 26'b01111100001100101101011110 :
  (x[23:13] == 1659) ? 26'b01111100000101100001101100 :
  (x[23:13] == 1660) ? 26'b01111011111110010110100110 :
  (x[23:13] == 1661) ? 26'b01111011110111001100010010 :
  (x[23:13] == 1662) ? 26'b01111011110000000010100110 :
  (x[23:13] == 1663) ? 26'b01111011101000111001100110 :
  (x[23:13] == 1664) ? 26'b01111011100001110001010000 :
  (x[23:13] == 1665) ? 26'b01111011011010101001101010 :
  (x[23:13] == 1666) ? 26'b01111011010011100010110000 :
  (x[23:13] == 1667) ? 26'b01111011001100011100100010 :
  (x[23:13] == 1668) ? 26'b01111011000101010110111000 :
  (x[23:13] == 1669) ? 26'b01111010111110010010000000 :
  (x[23:13] == 1670) ? 26'b01111010110111001101110010 :
  (x[23:13] == 1671) ? 26'b01111010110000001010001110 :
  (x[23:13] == 1672) ? 26'b01111010101001000111011000 :
  (x[23:13] == 1673) ? 26'b01111010100010000101001100 :
  (x[23:13] == 1674) ? 26'b01111010011011000011101100 :
  (x[23:13] == 1675) ? 26'b01111010010100000010110100 :
  (x[23:13] == 1676) ? 26'b01111010001101000010100100 :
  (x[23:13] == 1677) ? 26'b01111010000110000011000110 :
  (x[23:13] == 1678) ? 26'b01111001111111000100001100 :
  (x[23:13] == 1679) ? 26'b01111001111000000110000110 :
  (x[23:13] == 1680) ? 26'b01111001110001001000100000 :
  (x[23:13] == 1681) ? 26'b01111001101010001011101110 :
  (x[23:13] == 1682) ? 26'b01111001100011001111011110 :
  (x[23:13] == 1683) ? 26'b01111001011100010011111010 :
  (x[23:13] == 1684) ? 26'b01111001010101011001000110 :
  (x[23:13] == 1685) ? 26'b01111001001110011110110110 :
  (x[23:13] == 1686) ? 26'b01111001000111100101001110 :
  (x[23:13] == 1687) ? 26'b01111001000000101100010100 :
  (x[23:13] == 1688) ? 26'b01111000111001110100000110 :
  (x[23:13] == 1689) ? 26'b01111000110010111100011100 :
  (x[23:13] == 1690) ? 26'b01111000101100000101100100 :
  (x[23:13] == 1691) ? 26'b01111000100101001111001100 :
  (x[23:13] == 1692) ? 26'b01111000011110011001100000 :
  (x[23:13] == 1693) ? 26'b01111000010111100100100100 :
  (x[23:13] == 1694) ? 26'b01111000010000110000001010 :
  (x[23:13] == 1695) ? 26'b01111000001001111100011010 :
  (x[23:13] == 1696) ? 26'b01111000000011001001010100 :
  (x[23:13] == 1697) ? 26'b01110111111100010110111010 :
  (x[23:13] == 1698) ? 26'b01110111110101100101001000 :
  (x[23:13] == 1699) ? 26'b01110111101110110011111100 :
  (x[23:13] == 1700) ? 26'b01110111101000000011011000 :
  (x[23:13] == 1701) ? 26'b01110111100001010011011100 :
  (x[23:13] == 1702) ? 26'b01110111011010100100001010 :
  (x[23:13] == 1703) ? 26'b01110111010011110101100110 :
  (x[23:13] == 1704) ? 26'b01110111001101000111101000 :
  (x[23:13] == 1705) ? 26'b01110111000110011010010000 :
  (x[23:13] == 1706) ? 26'b01110110111111101101011100 :
  (x[23:13] == 1707) ? 26'b01110110111001000001011000 :
  (x[23:13] == 1708) ? 26'b01110110110010010101110110 :
  (x[23:13] == 1709) ? 26'b01110110101011101011000100 :
  (x[23:13] == 1710) ? 26'b01110110100101000000110110 :
  (x[23:13] == 1711) ? 26'b01110110011110010111001100 :
  (x[23:13] == 1712) ? 26'b01110110010111101110001010 :
  (x[23:13] == 1713) ? 26'b01110110010001000101110100 :
  (x[23:13] == 1714) ? 26'b01110110001010011110000100 :
  (x[23:13] == 1715) ? 26'b01110110000011110110111000 :
  (x[23:13] == 1716) ? 26'b01110101111101010000011000 :
  (x[23:13] == 1717) ? 26'b01110101110110101010011110 :
  (x[23:13] == 1718) ? 26'b01110101110000000101010000 :
  (x[23:13] == 1719) ? 26'b01110101101001100000100000 :
  (x[23:13] == 1720) ? 26'b01110101100010111100011100 :
  (x[23:13] == 1721) ? 26'b01110101011100011001000000 :
  (x[23:13] == 1722) ? 26'b01110101010101110110001100 :
  (x[23:13] == 1723) ? 26'b01110101001111010011111000 :
  (x[23:13] == 1724) ? 26'b01110101001000110010010000 :
  (x[23:13] == 1725) ? 26'b01110101000010010001010010 :
  (x[23:13] == 1726) ? 26'b01110100111011110000110100 :
  (x[23:13] == 1727) ? 26'b01110100110101010001000000 :
  (x[23:13] == 1728) ? 26'b01110100101110110001110000 :
  (x[23:13] == 1729) ? 26'b01110100101000010011001000 :
  (x[23:13] == 1730) ? 26'b01110100100001110101000010 :
  (x[23:13] == 1731) ? 26'b01110100011011010111101010 :
  (x[23:13] == 1732) ? 26'b01110100010100111010110100 :
  (x[23:13] == 1733) ? 26'b01110100001110011110100110 :
  (x[23:13] == 1734) ? 26'b01110100001000000011000010 :
  (x[23:13] == 1735) ? 26'b01110100000001100111111010 :
  (x[23:13] == 1736) ? 26'b01110011111011001101011100 :
  (x[23:13] == 1737) ? 26'b01110011110100110011100110 :
  (x[23:13] == 1738) ? 26'b01110011101110011010010100 :
  (x[23:13] == 1739) ? 26'b01110011101000000001101100 :
  (x[23:13] == 1740) ? 26'b01110011100001101001100000 :
  (x[23:13] == 1741) ? 26'b01110011011011010010000010 :
  (x[23:13] == 1742) ? 26'b01110011010100111011000110 :
  (x[23:13] == 1743) ? 26'b01110011001110100100101110 :
  (x[23:13] == 1744) ? 26'b01110011001000001110111110 :
  (x[23:13] == 1745) ? 26'b01110011000001111001110100 :
  (x[23:13] == 1746) ? 26'b01110010111011100101001010 :
  (x[23:13] == 1747) ? 26'b01110010110101010001001000 :
  (x[23:13] == 1748) ? 26'b01110010101110111101101110 :
  (x[23:13] == 1749) ? 26'b01110010101000101010110100 :
  (x[23:13] == 1750) ? 26'b01110010100010011000011110 :
  (x[23:13] == 1751) ? 26'b01110010011100000110110110 :
  (x[23:13] == 1752) ? 26'b01110010010101110101101000 :
  (x[23:13] == 1753) ? 26'b01110010001111100101000110 :
  (x[23:13] == 1754) ? 26'b01110010001001010101000110 :
  (x[23:13] == 1755) ? 26'b01110010000011000101101110 :
  (x[23:13] == 1756) ? 26'b01110001111100110110110100 :
  (x[23:13] == 1757) ? 26'b01110001110110101000100010 :
  (x[23:13] == 1758) ? 26'b01110001110000011010110000 :
  (x[23:13] == 1759) ? 26'b01110001101010001101100100 :
  (x[23:13] == 1760) ? 26'b01110001100100000000111110 :
  (x[23:13] == 1761) ? 26'b01110001011101110100111010 :
  (x[23:13] == 1762) ? 26'b01110001010111101001011100 :
  (x[23:13] == 1763) ? 26'b01110001010001011110100110 :
  (x[23:13] == 1764) ? 26'b01110001001011010100001110 :
  (x[23:13] == 1765) ? 26'b01110001000101001010010110 :
  (x[23:13] == 1766) ? 26'b01110000111111000001000100 :
  (x[23:13] == 1767) ? 26'b01110000111000111000011010 :
  (x[23:13] == 1768) ? 26'b01110000110010110000010110 :
  (x[23:13] == 1769) ? 26'b01110000101100101000110000 :
  (x[23:13] == 1770) ? 26'b01110000100110100001101110 :
  (x[23:13] == 1771) ? 26'b01110000100000011011001100 :
  (x[23:13] == 1772) ? 26'b01110000011010010101001110 :
  (x[23:13] == 1773) ? 26'b01110000010100001111111100 :
  (x[23:13] == 1774) ? 26'b01110000001110001011000010 :
  (x[23:13] == 1775) ? 26'b01110000001000000110110100 :
  (x[23:13] == 1776) ? 26'b01110000000010000011000100 :
  (x[23:13] == 1777) ? 26'b01101111111011111111111010 :
  (x[23:13] == 1778) ? 26'b01101111110101111101001110 :
  (x[23:13] == 1779) ? 26'b01101111101111111011001010 :
  (x[23:13] == 1780) ? 26'b01101111101001111001100010 :
  (x[23:13] == 1781) ? 26'b01101111100011111000100110 :
  (x[23:13] == 1782) ? 26'b01101111011101111000000100 :
  (x[23:13] == 1783) ? 26'b01101111010111111000001100 :
  (x[23:13] == 1784) ? 26'b01101111010001111000101110 :
  (x[23:13] == 1785) ? 26'b01101111001011111001110110 :
  (x[23:13] == 1786) ? 26'b01101111000101111011100000 :
  (x[23:13] == 1787) ? 26'b01101110111111111101110000 :
  (x[23:13] == 1788) ? 26'b01101110111010000000100100 :
  (x[23:13] == 1789) ? 26'b01101110110100000011110000 :
  (x[23:13] == 1790) ? 26'b01101110101110000111100000 :
  (x[23:13] == 1791) ? 26'b01101110101000001011111000 :
  (x[23:13] == 1792) ? 26'b01101110100010010000101110 :
  (x[23:13] == 1793) ? 26'b01101110011100010110001100 :
  (x[23:13] == 1794) ? 26'b01101110010110011100000110 :
  (x[23:13] == 1795) ? 26'b01101110010000100010011110 :
  (x[23:13] == 1796) ? 26'b01101110001010101001011100 :
  (x[23:13] == 1797) ? 26'b01101110000100110001000010 :
  (x[23:13] == 1798) ? 26'b01101101111110111001000100 :
  (x[23:13] == 1799) ? 26'b01101101111001000001100100 :
  (x[23:13] == 1800) ? 26'b01101101110011001010101010 :
  (x[23:13] == 1801) ? 26'b01101101101101010100001000 :
  (x[23:13] == 1802) ? 26'b01101101100111011110010000 :
  (x[23:13] == 1803) ? 26'b01101101100001101000111000 :
  (x[23:13] == 1804) ? 26'b01101101011011110100000110 :
  (x[23:13] == 1805) ? 26'b01101101010101111111101010 :
  (x[23:13] == 1806) ? 26'b01101101010000001011111010 :
  (x[23:13] == 1807) ? 26'b01101101001010011000100100 :
  (x[23:13] == 1808) ? 26'b01101101000100100101101110 :
  (x[23:13] == 1809) ? 26'b01101100111110110011011010 :
  (x[23:13] == 1810) ? 26'b01101100111001000001100110 :
  (x[23:13] == 1811) ? 26'b01101100110011010000010110 :
  (x[23:13] == 1812) ? 26'b01101100101101011111100110 :
  (x[23:13] == 1813) ? 26'b01101100100111101111011000 :
  (x[23:13] == 1814) ? 26'b01101100100001111111100100 :
  (x[23:13] == 1815) ? 26'b01101100011100010000011010 :
  (x[23:13] == 1816) ? 26'b01101100010110100001101000 :
  (x[23:13] == 1817) ? 26'b01101100010000110011011000 :
  (x[23:13] == 1818) ? 26'b01101100001011000101101010 :
  (x[23:13] == 1819) ? 26'b01101100000101011000011100 :
  (x[23:13] == 1820) ? 26'b01101011111111101011110000 :
  (x[23:13] == 1821) ? 26'b01101011111001111111100110 :
  (x[23:13] == 1822) ? 26'b01101011110100010011110100 :
  (x[23:13] == 1823) ? 26'b01101011101110101000100100 :
  (x[23:13] == 1824) ? 26'b01101011101000111101110100 :
  (x[23:13] == 1825) ? 26'b01101011100011010011100110 :
  (x[23:13] == 1826) ? 26'b01101011011101101001111000 :
  (x[23:13] == 1827) ? 26'b01101011011000000000101100 :
  (x[23:13] == 1828) ? 26'b01101011010010010111111010 :
  (x[23:13] == 1829) ? 26'b01101011001100101111101000 :
  (x[23:13] == 1830) ? 26'b01101011000111000111111000 :
  (x[23:13] == 1831) ? 26'b01101011000001100000101000 :
  (x[23:13] == 1832) ? 26'b01101010111011111001110110 :
  (x[23:13] == 1833) ? 26'b01101010110110010011100100 :
  (x[23:13] == 1834) ? 26'b01101010110000101101101110 :
  (x[23:13] == 1835) ? 26'b01101010101011001000100000 :
  (x[23:13] == 1836) ? 26'b01101010100101100011100100 :
  (x[23:13] == 1837) ? 26'b01101010011111111111010010 :
  (x[23:13] == 1838) ? 26'b01101010011010011011011000 :
  (x[23:13] == 1839) ? 26'b01101010010100111000000110 :
  (x[23:13] == 1840) ? 26'b01101010001111010101000110 :
  (x[23:13] == 1841) ? 26'b01101010001001110010101110 :
  (x[23:13] == 1842) ? 26'b01101010000100010000110100 :
  (x[23:13] == 1843) ? 26'b01101001111110101111011000 :
  (x[23:13] == 1844) ? 26'b01101001111001001110011000 :
  (x[23:13] == 1845) ? 26'b01101001110011101101111100 :
  (x[23:13] == 1846) ? 26'b01101001101110001101111000 :
  (x[23:13] == 1847) ? 26'b01101001101000101110011010 :
  (x[23:13] == 1848) ? 26'b01101001100011001111010100 :
  (x[23:13] == 1849) ? 26'b01101001011101110000101010 :
  (x[23:13] == 1850) ? 26'b01101001011000010010100110 :
  (x[23:13] == 1851) ? 26'b01101001010010110100111010 :
  (x[23:13] == 1852) ? 26'b01101001001101010111110010 :
  (x[23:13] == 1853) ? 26'b01101001000111111011000110 :
  (x[23:13] == 1854) ? 26'b01101001000010011110110100 :
  (x[23:13] == 1855) ? 26'b01101000111101000011000010 :
  (x[23:13] == 1856) ? 26'b01101000110111100111110000 :
  (x[23:13] == 1857) ? 26'b01101000110010001100111000 :
  (x[23:13] == 1858) ? 26'b01101000101100110010100110 :
  (x[23:13] == 1859) ? 26'b01101000100111011000101110 :
  (x[23:13] == 1860) ? 26'b01101000100001111111001110 :
  (x[23:13] == 1861) ? 26'b01101000011100100110010100 :
  (x[23:13] == 1862) ? 26'b01101000010111001101110100 :
  (x[23:13] == 1863) ? 26'b01101000010001110101101100 :
  (x[23:13] == 1864) ? 26'b01101000001100011110001100 :
  (x[23:13] == 1865) ? 26'b01101000000111000111000010 :
  (x[23:13] == 1866) ? 26'b01101000000001110000011010 :
  (x[23:13] == 1867) ? 26'b01100111111100011010001010 :
  (x[23:13] == 1868) ? 26'b01100111110111000100011000 :
  (x[23:13] == 1869) ? 26'b01100111110001101111001010 :
  (x[23:13] == 1870) ? 26'b01100111101100011010011000 :
  (x[23:13] == 1871) ? 26'b01100111100111000110000000 :
  (x[23:13] == 1872) ? 26'b01100111100001110010000110 :
  (x[23:13] == 1873) ? 26'b01100111011100011110100110 :
  (x[23:13] == 1874) ? 26'b01100111010111001011100100 :
  (x[23:13] == 1875) ? 26'b01100111010001111001000000 :
  (x[23:13] == 1876) ? 26'b01100111001100100110110110 :
  (x[23:13] == 1877) ? 26'b01100111000111010101001100 :
  (x[23:13] == 1878) ? 26'b01100111000010000100000000 :
  (x[23:13] == 1879) ? 26'b01100110111100110011001110 :
  (x[23:13] == 1880) ? 26'b01100110110111100010111010 :
  (x[23:13] == 1881) ? 26'b01100110110010010011001000 :
  (x[23:13] == 1882) ? 26'b01100110101101000011101100 :
  (x[23:13] == 1883) ? 26'b01100110100111110100101110 :
  (x[23:13] == 1884) ? 26'b01100110100010100110001000 :
  (x[23:13] == 1885) ? 26'b01100110011101011000000010 :
  (x[23:13] == 1886) ? 26'b01100110011000001010011100 :
  (x[23:13] == 1887) ? 26'b01100110010010111101001110 :
  (x[23:13] == 1888) ? 26'b01100110001101110000011110 :
  (x[23:13] == 1889) ? 26'b01100110001000100100000110 :
  (x[23:13] == 1890) ? 26'b01100110000011011000001110 :
  (x[23:13] == 1891) ? 26'b01100101111110001100110100 :
  (x[23:13] == 1892) ? 26'b01100101111001000001110010 :
  (x[23:13] == 1893) ? 26'b01100101110011110111001110 :
  (x[23:13] == 1894) ? 26'b01100101101110101101000110 :
  (x[23:13] == 1895) ? 26'b01100101101001100011011000 :
  (x[23:13] == 1896) ? 26'b01100101100100011010000100 :
  (x[23:13] == 1897) ? 26'b01100101011111010001010100 :
  (x[23:13] == 1898) ? 26'b01100101011010001000110110 :
  (x[23:13] == 1899) ? 26'b01100101010101000000111000 :
  (x[23:13] == 1900) ? 26'b01100101001111111001010110 :
  (x[23:13] == 1901) ? 26'b01100101001010110010001110 :
  (x[23:13] == 1902) ? 26'b01100101000101101011100100 :
  (x[23:13] == 1903) ? 26'b01100101000000100101011000 :
  (x[23:13] == 1904) ? 26'b01100100111011011111100100 :
  (x[23:13] == 1905) ? 26'b01100100110110011010000110 :
  (x[23:13] == 1906) ? 26'b01100100110001010101001000 :
  (x[23:13] == 1907) ? 26'b01100100101100010000101010 :
  (x[23:13] == 1908) ? 26'b01100100100111001100100000 :
  (x[23:13] == 1909) ? 26'b01100100100010001000111000 :
  (x[23:13] == 1910) ? 26'b01100100011101000101100110 :
  (x[23:13] == 1911) ? 26'b01100100011000000010110010 :
  (x[23:13] == 1912) ? 26'b01100100010011000000010100 :
  (x[23:13] == 1913) ? 26'b01100100001101111110010110 :
  (x[23:13] == 1914) ? 26'b01100100001000111100110000 :
  (x[23:13] == 1915) ? 26'b01100100000011111011101000 :
  (x[23:13] == 1916) ? 26'b01100011111110111010111000 :
  (x[23:13] == 1917) ? 26'b01100011111001111010100010 :
  (x[23:13] == 1918) ? 26'b01100011110100111010100110 :
  (x[23:13] == 1919) ? 26'b01100011101111111011001000 :
  (x[23:13] == 1920) ? 26'b01100011101010111100000100 :
  (x[23:13] == 1921) ? 26'b01100011100101111101011100 :
  (x[23:13] == 1922) ? 26'b01100011100000111111001010 :
  (x[23:13] == 1923) ? 26'b01100011011100000001010110 :
  (x[23:13] == 1924) ? 26'b01100011010111000011111010 :
  (x[23:13] == 1925) ? 26'b01100011010010000110111010 :
  (x[23:13] == 1926) ? 26'b01100011001101001010010010 :
  (x[23:13] == 1927) ? 26'b01100011001000001110001010 :
  (x[23:13] == 1928) ? 26'b01100011000011010010010110 :
  (x[23:13] == 1929) ? 26'b01100010111110010110111110 :
  (x[23:13] == 1930) ? 26'b01100010111001011011111110 :
  (x[23:13] == 1931) ? 26'b01100010110100100001100000 :
  (x[23:13] == 1932) ? 26'b01100010101111100111010110 :
  (x[23:13] == 1933) ? 26'b01100010101010101101100110 :
  (x[23:13] == 1934) ? 26'b01100010100101110100010010 :
  (x[23:13] == 1935) ? 26'b01100010100000111011011010 :
  (x[23:13] == 1936) ? 26'b01100010011100000010110110 :
  (x[23:13] == 1937) ? 26'b01100010010111001010110010 :
  (x[23:13] == 1938) ? 26'b01100010010010010011000000 :
  (x[23:13] == 1939) ? 26'b01100010001101011011101100 :
  (x[23:13] == 1940) ? 26'b01100010001000100100110100 :
  (x[23:13] == 1941) ? 26'b01100010000011101110010100 :
  (x[23:13] == 1942) ? 26'b01100001111110111000001100 :
  (x[23:13] == 1943) ? 26'b01100001111010000010011110 :
  (x[23:13] == 1944) ? 26'b01100001110101001101001010 :
  (x[23:13] == 1945) ? 26'b01100001110000011000010000 :
  (x[23:13] == 1946) ? 26'b01100001101011100011110010 :
  (x[23:13] == 1947) ? 26'b01100001100110101111100110 :
  (x[23:13] == 1948) ? 26'b01100001100001111011111000 :
  (x[23:13] == 1949) ? 26'b01100001011101001000100010 :
  (x[23:13] == 1950) ? 26'b01100001011000010101100110 :
  (x[23:13] == 1951) ? 26'b01100001010011100011000100 :
  (x[23:13] == 1952) ? 26'b01100001001110110000110110 :
  (x[23:13] == 1953) ? 26'b01100001001001111111001000 :
  (x[23:13] == 1954) ? 26'b01100001000101001101110000 :
  (x[23:13] == 1955) ? 26'b01100001000000011100110010 :
  (x[23:13] == 1956) ? 26'b01100000111011101100001100 :
  (x[23:13] == 1957) ? 26'b01100000110110111011111110 :
  (x[23:13] == 1958) ? 26'b01100000110010001100001100 :
  (x[23:13] == 1959) ? 26'b01100000101101011100101110 :
  (x[23:13] == 1960) ? 26'b01100000101000101101101000 :
  (x[23:13] == 1961) ? 26'b01100000100011111111000000 :
  (x[23:13] == 1962) ? 26'b01100000011111010000101110 :
  (x[23:13] == 1963) ? 26'b01100000011010100010111000 :
  (x[23:13] == 1964) ? 26'b01100000010101110101011010 :
  (x[23:13] == 1965) ? 26'b01100000010001001000010000 :
  (x[23:13] == 1966) ? 26'b01100000001100011011100100 :
  (x[23:13] == 1967) ? 26'b01100000000111101111001100 :
  (x[23:13] == 1968) ? 26'b01100000000011000011001100 :
  (x[23:13] == 1969) ? 26'b01011111111110010111101000 :
  (x[23:13] == 1970) ? 26'b01011111111001101100011110 :
  (x[23:13] == 1971) ? 26'b01011111110101000001100110 :
  (x[23:13] == 1972) ? 26'b01011111110000010111001100 :
  (x[23:13] == 1973) ? 26'b01011111101011101101000110 :
  (x[23:13] == 1974) ? 26'b01011111100111000011011000 :
  (x[23:13] == 1975) ? 26'b01011111100010011010000000 :
  (x[23:13] == 1976) ? 26'b01011111011101110001000100 :
  (x[23:13] == 1977) ? 26'b01011111011001001000100010 :
  (x[23:13] == 1978) ? 26'b01011111010100100000010010 :
  (x[23:13] == 1979) ? 26'b01011111001111111000100000 :
  (x[23:13] == 1980) ? 26'b01011111001011010001000010 :
  (x[23:13] == 1981) ? 26'b01011111000110101001111110 :
  (x[23:13] == 1982) ? 26'b01011111000010000011010010 :
  (x[23:13] == 1983) ? 26'b01011110111101011100111110 :
  (x[23:13] == 1984) ? 26'b01011110111000110110111110 :
  (x[23:13] == 1985) ? 26'b01011110110100010001011000 :
  (x[23:13] == 1986) ? 26'b01011110101111101100001100 :
  (x[23:13] == 1987) ? 26'b01011110101011000111010100 :
  (x[23:13] == 1988) ? 26'b01011110100110100010111000 :
  (x[23:13] == 1989) ? 26'b01011110100001111110110000 :
  (x[23:13] == 1990) ? 26'b01011110011101011011000000 :
  (x[23:13] == 1991) ? 26'b01011110011000110111100100 :
  (x[23:13] == 1992) ? 26'b01011110010100010100100110 :
  (x[23:13] == 1993) ? 26'b01011110001111110001111100 :
  (x[23:13] == 1994) ? 26'b01011110001011001111101010 :
  (x[23:13] == 1995) ? 26'b01011110000110101101110000 :
  (x[23:13] == 1996) ? 26'b01011110000010001100001110 :
  (x[23:13] == 1997) ? 26'b01011101111101101011000000 :
  (x[23:13] == 1998) ? 26'b01011101111001001010001010 :
  (x[23:13] == 1999) ? 26'b01011101110100101001101000 :
  (x[23:13] == 2000) ? 26'b01011101110000001001100000 :
  (x[23:13] == 2001) ? 26'b01011101101011101001110010 :
  (x[23:13] == 2002) ? 26'b01011101100111001010011010 :
  (x[23:13] == 2003) ? 26'b01011101100010101011010100 :
  (x[23:13] == 2004) ? 26'b01011101011110001100101100 :
  (x[23:13] == 2005) ? 26'b01011101011001101110010110 :
  (x[23:13] == 2006) ? 26'b01011101010101010000011000 :
  (x[23:13] == 2007) ? 26'b01011101010000110010110100 :
  (x[23:13] == 2008) ? 26'b01011101001100010101011110 :
  (x[23:13] == 2009) ? 26'b01011101000111111000100110 :
  (x[23:13] == 2010) ? 26'b01011101000011011100000010 :
  (x[23:13] == 2011) ? 26'b01011100111110111111111010 :
  (x[23:13] == 2012) ? 26'b01011100111010100100000000 :
  (x[23:13] == 2013) ? 26'b01011100110110001000100010 :
  (x[23:13] == 2014) ? 26'b01011100110001101101011000 :
  (x[23:13] == 2015) ? 26'b01011100101101010010101100 :
  (x[23:13] == 2016) ? 26'b01011100101000111000001100 :
  (x[23:13] == 2017) ? 26'b01011100100100011110001010 :
  (x[23:13] == 2018) ? 26'b01011100100000000100011110 :
  (x[23:13] == 2019) ? 26'b01011100011011101011000010 :
  (x[23:13] == 2020) ? 26'b01011100010111010001111110 :
  (x[23:13] == 2021) ? 26'b01011100010010111001001110 :
  (x[23:13] == 2022) ? 26'b01011100001110100000111100 :
  (x[23:13] == 2023) ? 26'b01011100001010001000111100 :
  (x[23:13] == 2024) ? 26'b01011100000101110001010010 :
  (x[23:13] == 2025) ? 26'b01011100000001011010000000 :
  (x[23:13] == 2026) ? 26'b01011011111101000011000000 :
  (x[23:13] == 2027) ? 26'b01011011111000101100011010 :
  (x[23:13] == 2028) ? 26'b01011011110100010110001010 :
  (x[23:13] == 2029) ? 26'b01011011110000000000001110 :
  (x[23:13] == 2030) ? 26'b01011011101011101010101000 :
  (x[23:13] == 2031) ? 26'b01011011100111010101011000 :
  (x[23:13] == 2032) ? 26'b01011011100011000000011100 :
  (x[23:13] == 2033) ? 26'b01011011011110101011111000 :
  (x[23:13] == 2034) ? 26'b01011011011010010111101100 :
  (x[23:13] == 2035) ? 26'b01011011010110000011110110 :
  (x[23:13] == 2036) ? 26'b01011011010001110000010000 :
  (x[23:13] == 2037) ? 26'b01011011001101011101000100 :
  (x[23:13] == 2038) ? 26'b01011011001001001010001010 :
  (x[23:13] == 2039) ? 26'b01011011000100110111101000 :
  (x[23:13] == 2040) ? 26'b01011011000000100101011000 :
  (x[23:13] == 2041) ? 26'b01011010111100010011100100 :
  (x[23:13] == 2042) ? 26'b01011010111000000010000100 :
  (x[23:13] == 2043) ? 26'b01011010110011110000110100 :
  (x[23:13] == 2044) ? 26'b01011010101111011111111100 :
  (x[23:13] == 2045) ? 26'b01011010101011001111100000 :
  (x[23:13] == 2046) ? 26'b01011010100110111111010000 :
  26'b01011010100010101111011100 ;
  
  
 
  wire state;
  assign state = x[23]; //1ならodd,0ならeven
  
  wire [25:0] manx;
  assign manx = {3'b001, mx};


//小数点は23*2より、下から47bit目と46bit目の境目。
//偶数(つまり指数部の最下位が0)の時は、割る4ゆえ49と48の境目になり、
//奇数(つまり指数部の最下位が1)の時は、割る8ゆえ50と49の境目になる.
  wire [50:0] b;
  assign b = manx * cube_reg;
  

//小数点は上位2bit目と3bit目との間。結果は、01.hogeとなっているはず      
  wire [25:0] m_gap;
  assign m_gap = state ? three_reg - b[50:25]  : three_reg - b[49:24] ;  //bの下位1bitは捨てうる  
  wire [22:0] my;
  assign my = m_gap[23:1];
  
  wire [7:0] eodd;
  assign eodd = 8'd255 - ex[7:0];
  wire [7:0] ey;
  assign ey = state ? (8'd62 + {1'b0, eodd[7:1]}) : (8'd190 - {1'b0, ex[7:1]}) ;  

  wire [31:0] x_sqrt_inv;
  assign x_sqrt_inv = {sx, ey, my};

  logic [31:0] tmp;
  
// x*x^(-1/2)=x^1/2　　
  fmul u1(x, tmp, y);

always @(posedge clk) begin
    three_reg <= three;
    cube_reg <= cube;
    tmp <= x_sqrt_inv;
end
  
endmodule
