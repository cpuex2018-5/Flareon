`timescale 1ns / 1ps

//とりあえず組み合わせ回路で実現しようか

module finv(
  input clk,
  input wire [31:0] x,
  output wire [31:0] y);
  
  wire sx;
  wire [7:0] ex;
  wire [22:0] mx;
  
  assign {sx,ex,mx}=x;
  
  //25bit_verに対応させた
  wire [24:0] twice;
  wire [24:0] square;

  logic [24:0] twice_table [0:2047]; 
  logic [24:0] square_table [0:2047];
  
  //テーブルをもとに作成
  initial begin
      twice_table[0] = 25'b1111111111110000000000010;
      twice_table[1] = 25'b1111111111010000000010010;
      twice_table[2] = 25'b1111111110110000000110010;
      twice_table[3] = 25'b1111111110010000001100010;
      twice_table[4] = 25'b1111111101110000010100010;
      twice_table[5] = 25'b1111111101010000011110010;
      twice_table[6] = 25'b1111111100110000101010000;
      twice_table[7] = 25'b1111111100010000111000000;
      twice_table[8] = 25'b1111111011110001001000000;
      twice_table[9] = 25'b1111111011010001011001110;
      twice_table[10] = 25'b1111111010110001101101110;
      twice_table[11] = 25'b1111111010010010000011100;
      twice_table[12] = 25'b1111111001110010011011010;
      twice_table[13] = 25'b1111111001010010110101000;
      twice_table[14] = 25'b1111111000110011010000110;
      twice_table[15] = 25'b1111111000010011101110100;
      twice_table[16] = 25'b1111110111110100001110000;
      twice_table[17] = 25'b1111110111010100101111110;
      twice_table[18] = 25'b1111110110110101010011010;
      twice_table[19] = 25'b1111110110010101111000110;
      twice_table[20] = 25'b1111110101110110100000000;
      twice_table[21] = 25'b1111110101010111001001100;
      twice_table[22] = 25'b1111110100110111110100110;
      twice_table[23] = 25'b1111110100011000100010000;
      twice_table[24] = 25'b1111110011111001010001010;
      twice_table[25] = 25'b1111110011011010000010010;
      twice_table[26] = 25'b1111110010111010110101010;
      twice_table[27] = 25'b1111110010011011101010010;
      twice_table[28] = 25'b1111110001111100100001000;
      twice_table[29] = 25'b1111110001011101011010000;
      twice_table[30] = 25'b1111110000111110010100100;
      twice_table[31] = 25'b1111110000011111010001010;
      twice_table[32] = 25'b1111110000000000001111110;
      twice_table[33] = 25'b1111101111100001010000010;
      twice_table[34] = 25'b1111101111000010010010100;
      twice_table[35] = 25'b1111101110100011010110110;
      twice_table[36] = 25'b1111101110000100011101000;
      twice_table[37] = 25'b1111101101100101100101000;
      twice_table[38] = 25'b1111101101000110101111000;
      twice_table[39] = 25'b1111101100100111111010110;
      twice_table[40] = 25'b1111101100001001001000100;
      twice_table[41] = 25'b1111101011101010011000000;
      twice_table[42] = 25'b1111101011001011101001100;
      twice_table[43] = 25'b1111101010101100111101000;
      twice_table[44] = 25'b1111101010001110010010010;
      twice_table[45] = 25'b1111101001101111101001010;
      twice_table[46] = 25'b1111101001010001000010010;
      twice_table[47] = 25'b1111101000110010011101000;
      twice_table[48] = 25'b1111101000010011111001110;
      twice_table[49] = 25'b1111100111110101011000100;
      twice_table[50] = 25'b1111100111010110111001000;
      twice_table[51] = 25'b1111100110111000011011010;
      twice_table[52] = 25'b1111100110011001111111010;
      twice_table[53] = 25'b1111100101111011100101100;
      twice_table[54] = 25'b1111100101011101001101010;
      twice_table[55] = 25'b1111100100111110110111000;
      twice_table[56] = 25'b1111100100100000100010100;
      twice_table[57] = 25'b1111100100000010010000000;
      twice_table[58] = 25'b1111100011100011111111010;
      twice_table[59] = 25'b1111100011000101110000010;
      twice_table[60] = 25'b1111100010100111100011010;
      twice_table[61] = 25'b1111100010001001011000000;
      twice_table[62] = 25'b1111100001101011001110100;
      twice_table[63] = 25'b1111100001001101000111000;
      twice_table[64] = 25'b1111100000101111000001010;
      twice_table[65] = 25'b1111100000010000111101010;
      twice_table[66] = 25'b1111011111110010111011010;
      twice_table[67] = 25'b1111011111010100111010110;
      twice_table[68] = 25'b1111011110110110111100100;
      twice_table[69] = 25'b1111011110011000111111110;
      twice_table[70] = 25'b1111011101111011000100110;
      twice_table[71] = 25'b1111011101011101001011110;
      twice_table[72] = 25'b1111011100111111010100100;
      twice_table[73] = 25'b1111011100100001011111000;
      twice_table[74] = 25'b1111011100000011101011100;
      twice_table[75] = 25'b1111011011100101111001100;
      twice_table[76] = 25'b1111011011001000001001100;
      twice_table[77] = 25'b1111011010101010011011010;
      twice_table[78] = 25'b1111011010001100101110110;
      twice_table[79] = 25'b1111011001101111000100000;
      twice_table[80] = 25'b1111011001010001011011010;
      twice_table[81] = 25'b1111011000110011110100000;
      twice_table[82] = 25'b1111011000010110001110110;
      twice_table[83] = 25'b1111010111111000101011000;
      twice_table[84] = 25'b1111010111011011001001010;
      twice_table[85] = 25'b1111010110111101101001010;
      twice_table[86] = 25'b1111010110100000001011000;
      twice_table[87] = 25'b1111010110000010101110100;
      twice_table[88] = 25'b1111010101100101010011110;
      twice_table[89] = 25'b1111010101000111111010110;
      twice_table[90] = 25'b1111010100101010100011110;
      twice_table[91] = 25'b1111010100001101001110010;
      twice_table[92] = 25'b1111010011101111111010100;
      twice_table[93] = 25'b1111010011010010101000100;
      twice_table[94] = 25'b1111010010110101011000010;
      twice_table[95] = 25'b1111010010011000001010000;
      twice_table[96] = 25'b1111010001111010111101010;
      twice_table[97] = 25'b1111010001011101110010010;
      twice_table[98] = 25'b1111010001000000101001000;
      twice_table[99] = 25'b1111010000100011100001100;
      twice_table[100] = 25'b1111010000000110011011110;
      twice_table[101] = 25'b1111001111101001010111110;
      twice_table[102] = 25'b1111001111001100010101100;
      twice_table[103] = 25'b1111001110101111010101000;
      twice_table[104] = 25'b1111001110010010010110000;
      twice_table[105] = 25'b1111001101110101011001000;
      twice_table[106] = 25'b1111001101011000011101100;
      twice_table[107] = 25'b1111001100111011100100000;
      twice_table[108] = 25'b1111001100011110101100000;
      twice_table[109] = 25'b1111001100000001110101110;
      twice_table[110] = 25'b1111001011100101000001010;
      twice_table[111] = 25'b1111001011001000001110010;
      twice_table[112] = 25'b1111001010101011011101010;
      twice_table[113] = 25'b1111001010001110101101110;
      twice_table[114] = 25'b1111001001110010000000000;
      twice_table[115] = 25'b1111001001010101010100000;
      twice_table[116] = 25'b1111001000111000101001110;
      twice_table[117] = 25'b1111001000011100000001000;
      twice_table[118] = 25'b1111000111111111011010010;
      twice_table[119] = 25'b1111000111100010110101000;
      twice_table[120] = 25'b1111000111000110010001100;
      twice_table[121] = 25'b1111000110101001101111100;
      twice_table[122] = 25'b1111000110001101001111010;
      twice_table[123] = 25'b1111000101110000110000110;
      twice_table[124] = 25'b1111000101010100010100000;
      twice_table[125] = 25'b1111000100110111111000110;
      twice_table[126] = 25'b1111000100011011011111010;
      twice_table[127] = 25'b1111000011111111000111100;
      twice_table[128] = 25'b1111000011100010110001010;
      twice_table[129] = 25'b1111000011000110011101000;
      twice_table[130] = 25'b1111000010101010001010000;
      twice_table[131] = 25'b1111000010001101111001000;
      twice_table[132] = 25'b1111000001110001101001100;
      twice_table[133] = 25'b1111000001010101011011100;
      twice_table[134] = 25'b1111000000111001001111100;
      twice_table[135] = 25'b1111000000011101000101000;
      twice_table[136] = 25'b1111000000000000111100000;
      twice_table[137] = 25'b1110111111100100110100110;
      twice_table[138] = 25'b1110111111001000101111010;
      twice_table[139] = 25'b1110111110101100101011010;
      twice_table[140] = 25'b1110111110010000101001000;
      twice_table[141] = 25'b1110111101110100101000010;
      twice_table[142] = 25'b1110111101011000101001010;
      twice_table[143] = 25'b1110111100111100101011110;
      twice_table[144] = 25'b1110111100100000110000000;
      twice_table[145] = 25'b1110111100000100110110000;
      twice_table[146] = 25'b1110111011101000111101100;
      twice_table[147] = 25'b1110111011001101000110100;
      twice_table[148] = 25'b1110111010110001010001010;
      twice_table[149] = 25'b1110111010010101011101110;
      twice_table[150] = 25'b1110111001111001101011110;
      twice_table[151] = 25'b1110111001011101111011010;
      twice_table[152] = 25'b1110111001000010001100100;
      twice_table[153] = 25'b1110111000100110011111010;
      twice_table[154] = 25'b1110111000001010110011110;
      twice_table[155] = 25'b1110110111101111001001110;
      twice_table[156] = 25'b1110110111010011100001100;
      twice_table[157] = 25'b1110110110110111111010110;
      twice_table[158] = 25'b1110110110011100010101110;
      twice_table[159] = 25'b1110110110000000110010000;
      twice_table[160] = 25'b1110110101100101010000010;
      twice_table[161] = 25'b1110110101001001101111110;
      twice_table[162] = 25'b1110110100101110010001000;
      twice_table[163] = 25'b1110110100010010110100000;
      twice_table[164] = 25'b1110110011110111011000010;
      twice_table[165] = 25'b1110110011011011111110010;
      twice_table[166] = 25'b1110110011000000100110000;
      twice_table[167] = 25'b1110110010100101001111000;
      twice_table[168] = 25'b1110110010001001111001110;
      twice_table[169] = 25'b1110110001101110100110010;
      twice_table[170] = 25'b1110110001010011010100000;
      twice_table[171] = 25'b1110110000111000000011100;
      twice_table[172] = 25'b1110110000011100110100110;
      twice_table[173] = 25'b1110110000000001100111010;
      twice_table[174] = 25'b1110101111100110011011100;
      twice_table[175] = 25'b1110101111001011010001010;
      twice_table[176] = 25'b1110101110110000001000100;
      twice_table[177] = 25'b1110101110010101000001100;
      twice_table[178] = 25'b1110101101111001111011110;
      twice_table[179] = 25'b1110101101011110110111110;
      twice_table[180] = 25'b1110101101000011110101010;
      twice_table[181] = 25'b1110101100101000110100100;
      twice_table[182] = 25'b1110101100001101110101010;
      twice_table[183] = 25'b1110101011110010110111010;
      twice_table[184] = 25'b1110101011010111111011000;
      twice_table[185] = 25'b1110101010111101000000010;
      twice_table[186] = 25'b1110101010100010000111010;
      twice_table[187] = 25'b1110101010000111001111100;
      twice_table[188] = 25'b1110101001101100011001100;
      twice_table[189] = 25'b1110101001010001100101000;
      twice_table[190] = 25'b1110101000110110110010000;
      twice_table[191] = 25'b1110101000011100000000100;
      twice_table[192] = 25'b1110101000000001010000100;
      twice_table[193] = 25'b1110100111100110100010000;
      twice_table[194] = 25'b1110100111001011110101000;
      twice_table[195] = 25'b1110100110110001001001110;
      twice_table[196] = 25'b1110100110010110011111110;
      twice_table[197] = 25'b1110100101111011110111100;
      twice_table[198] = 25'b1110100101100001010000110;
      twice_table[199] = 25'b1110100101000110101011010;
      twice_table[200] = 25'b1110100100101100000111100;
      twice_table[201] = 25'b1110100100010001100101010;
      twice_table[202] = 25'b1110100011110111000100100;
      twice_table[203] = 25'b1110100011011100100101010;
      twice_table[204] = 25'b1110100011000010000111100;
      twice_table[205] = 25'b1110100010100111101011010;
      twice_table[206] = 25'b1110100010001101010000100;
      twice_table[207] = 25'b1110100001110010110111010;
      twice_table[208] = 25'b1110100001011000011111100;
      twice_table[209] = 25'b1110100000111110001001010;
      twice_table[210] = 25'b1110100000100011110100100;
      twice_table[211] = 25'b1110100000001001100001000;
      twice_table[212] = 25'b1110011111101111001111010;
      twice_table[213] = 25'b1110011111010100111111000;
      twice_table[214] = 25'b1110011110111010110000010;
      twice_table[215] = 25'b1110011110100000100010110;
      twice_table[216] = 25'b1110011110000110010111000;
      twice_table[217] = 25'b1110011101101100001100100;
      twice_table[218] = 25'b1110011101010010000011110;
      twice_table[219] = 25'b1110011100110111111100010;
      twice_table[220] = 25'b1110011100011101110110010;
      twice_table[221] = 25'b1110011100000011110001110;
      twice_table[222] = 25'b1110011011101001101110110;
      twice_table[223] = 25'b1110011011001111101101010;
      twice_table[224] = 25'b1110011010110101101101010;
      twice_table[225] = 25'b1110011010011011101110100;
      twice_table[226] = 25'b1110011010000001110001100;
      twice_table[227] = 25'b1110011001100111110101110;
      twice_table[228] = 25'b1110011001001101111011100;
      twice_table[229] = 25'b1110011000110100000010110;
      twice_table[230] = 25'b1110011000011010001011100;
      twice_table[231] = 25'b1110011000000000010101100;
      twice_table[232] = 25'b1110010111100110100001010;
      twice_table[233] = 25'b1110010111001100101110010;
      twice_table[234] = 25'b1110010110110010111100110;
      twice_table[235] = 25'b1110010110011001001100100;
      twice_table[236] = 25'b1110010101111111011110000;
      twice_table[237] = 25'b1110010101100101110000110;
      twice_table[238] = 25'b1110010101001100000101000;
      twice_table[239] = 25'b1110010100110010011010110;
      twice_table[240] = 25'b1110010100011000110001110;
      twice_table[241] = 25'b1110010011111111001010010;
      twice_table[242] = 25'b1110010011100101100100010;
      twice_table[243] = 25'b1110010011001011111111110;
      twice_table[244] = 25'b1110010010110010011100100;
      twice_table[245] = 25'b1110010010011000111010110;
      twice_table[246] = 25'b1110010001111111011010100;
      twice_table[247] = 25'b1110010001100101111011100;
      twice_table[248] = 25'b1110010001001100011110010;
      twice_table[249] = 25'b1110010000110011000010000;
      twice_table[250] = 25'b1110010000011001100111100;
      twice_table[251] = 25'b1110010000000000001110010;
      twice_table[252] = 25'b1110001111100110110110100;
      twice_table[253] = 25'b1110001111001101100000000;
      twice_table[254] = 25'b1110001110110100001011000;
      twice_table[255] = 25'b1110001110011010110111100;
      twice_table[256] = 25'b1110001110000001100101010;
      twice_table[257] = 25'b1110001101101000010100100;
      twice_table[258] = 25'b1110001101001111000101010;
      twice_table[259] = 25'b1110001100110101110111010;
      twice_table[260] = 25'b1110001100011100101010110;
      twice_table[261] = 25'b1110001100000011011111100;
      twice_table[262] = 25'b1110001011101010010101110;
      twice_table[263] = 25'b1110001011010001001101010;
      twice_table[264] = 25'b1110001010111000000110010;
      twice_table[265] = 25'b1110001010011111000000110;
      twice_table[266] = 25'b1110001010000101111100100;
      twice_table[267] = 25'b1110001001101100111001110;
      twice_table[268] = 25'b1110001001010011111000010;
      twice_table[269] = 25'b1110001000111010111000010;
      twice_table[270] = 25'b1110001000100001111001100;
      twice_table[271] = 25'b1110001000001000111100010;
      twice_table[272] = 25'b1110000111110000000000010;
      twice_table[273] = 25'b1110000111010111000101110;
      twice_table[274] = 25'b1110000110111110001100100;
      twice_table[275] = 25'b1110000110100101010100110;
      twice_table[276] = 25'b1110000110001100011110010;
      twice_table[277] = 25'b1110000101110011101001010;
      twice_table[278] = 25'b1110000101011010110101100;
      twice_table[279] = 25'b1110000101000010000011000;
      twice_table[280] = 25'b1110000100101001010010010;
      twice_table[281] = 25'b1110000100010000100010100;
      twice_table[282] = 25'b1110000011110111110100010;
      twice_table[283] = 25'b1110000011011111000111010;
      twice_table[284] = 25'b1110000011000110011011110;
      twice_table[285] = 25'b1110000010101101110001100;
      twice_table[286] = 25'b1110000010010101001000110;
      twice_table[287] = 25'b1110000001111100100001010;
      twice_table[288] = 25'b1110000001100011111011000;
      twice_table[289] = 25'b1110000001001011010110010;
      twice_table[290] = 25'b1110000000110010110011000;
      twice_table[291] = 25'b1110000000011010010000110;
      twice_table[292] = 25'b1110000000000001110000000;
      twice_table[293] = 25'b1101111111101001010000100;
      twice_table[294] = 25'b1101111111010000110010100;
      twice_table[295] = 25'b1101111110111000010101110;
      twice_table[296] = 25'b1101111110011111111010010;
      twice_table[297] = 25'b1101111110000111100000010;
      twice_table[298] = 25'b1101111101101111000111100;
      twice_table[299] = 25'b1101111101010110110000000;
      twice_table[300] = 25'b1101111100111110011010000;
      twice_table[301] = 25'b1101111100100110000101010;
      twice_table[302] = 25'b1101111100001101110001110;
      twice_table[303] = 25'b1101111011110101011111110;
      twice_table[304] = 25'b1101111011011101001110110;
      twice_table[305] = 25'b1101111011000100111111010;
      twice_table[306] = 25'b1101111010101100110001010;
      twice_table[307] = 25'b1101111010010100100100010;
      twice_table[308] = 25'b1101111001111100011000110;
      twice_table[309] = 25'b1101111001100100001110100;
      twice_table[310] = 25'b1101111001001100000101110;
      twice_table[311] = 25'b1101111000110011111110000;
      twice_table[312] = 25'b1101111000011011110111110;
      twice_table[313] = 25'b1101111000000011110010110;
      twice_table[314] = 25'b1101110111101011101111010;
      twice_table[315] = 25'b1101110111010011101100110;
      twice_table[316] = 25'b1101110110111011101011110;
      twice_table[317] = 25'b1101110110100011101100000;
      twice_table[318] = 25'b1101110110001011101101100;
      twice_table[319] = 25'b1101110101110011110000010;
      twice_table[320] = 25'b1101110101011011110100100;
      twice_table[321] = 25'b1101110101000011111001110;
      twice_table[322] = 25'b1101110100101100000000100;
      twice_table[323] = 25'b1101110100010100001000100;
      twice_table[324] = 25'b1101110011111100010001110;
      twice_table[325] = 25'b1101110011100100011100010;
      twice_table[326] = 25'b1101110011001100101000010;
      twice_table[327] = 25'b1101110010110100110101010;
      twice_table[328] = 25'b1101110010011101000011110;
      twice_table[329] = 25'b1101110010000101010011100;
      twice_table[330] = 25'b1101110001101101100100010;
      twice_table[331] = 25'b1101110001010101110110100;
      twice_table[332] = 25'b1101110000111110001010010;
      twice_table[333] = 25'b1101110000100110011111000;
      twice_table[334] = 25'b1101110000001110110101000;
      twice_table[335] = 25'b1101101111110111001100010;
      twice_table[336] = 25'b1101101111011111100101000;
      twice_table[337] = 25'b1101101111000111111110110;
      twice_table[338] = 25'b1101101110110000011010000;
      twice_table[339] = 25'b1101101110011000110110010;
      twice_table[340] = 25'b1101101110000001010100000;
      twice_table[341] = 25'b1101101101101001110011000;
      twice_table[342] = 25'b1101101101010010010011010;
      twice_table[343] = 25'b1101101100111010110100100;
      twice_table[344] = 25'b1101101100100011010111010;
      twice_table[345] = 25'b1101101100001011111011010;
      twice_table[346] = 25'b1101101011110100100000100;
      twice_table[347] = 25'b1101101011011101000111000;
      twice_table[348] = 25'b1101101011000101101110100;
      twice_table[349] = 25'b1101101010101110010111100;
      twice_table[350] = 25'b1101101010010111000001110;
      twice_table[351] = 25'b1101101001111111101101010;
      twice_table[352] = 25'b1101101001101000011010000;
      twice_table[353] = 25'b1101101001010001000111110;
      twice_table[354] = 25'b1101101000111001110111000;
      twice_table[355] = 25'b1101101000100010100111100;
      twice_table[356] = 25'b1101101000001011011001000;
      twice_table[357] = 25'b1101100111110100001100000;
      twice_table[358] = 25'b1101100111011101000000000;
      twice_table[359] = 25'b1101100111000101110101100;
      twice_table[360] = 25'b1101100110101110101100000;
      twice_table[361] = 25'b1101100110010111100011110;
      twice_table[362] = 25'b1101100110000000011101000;
      twice_table[363] = 25'b1101100101101001010111010;
      twice_table[364] = 25'b1101100101010010010010110;
      twice_table[365] = 25'b1101100100111011001111010;
      twice_table[366] = 25'b1101100100100100001101010;
      twice_table[367] = 25'b1101100100001101001100100;
      twice_table[368] = 25'b1101100011110110001100110;
      twice_table[369] = 25'b1101100011011111001110100;
      twice_table[370] = 25'b1101100011001000010001010;
      twice_table[371] = 25'b1101100010110001010101010;
      twice_table[372] = 25'b1101100010011010011010100;
      twice_table[373] = 25'b1101100010000011100001000;
      twice_table[374] = 25'b1101100001101100101000110;
      twice_table[375] = 25'b1101100001010101110001100;
      twice_table[376] = 25'b1101100000111110111011100;
      twice_table[377] = 25'b1101100000101000000110110;
      twice_table[378] = 25'b1101100000010001010011010;
      twice_table[379] = 25'b1101011111111010100001000;
      twice_table[380] = 25'b1101011111100011110000000;
      twice_table[381] = 25'b1101011111001101000000000;
      twice_table[382] = 25'b1101011110110110010001010;
      twice_table[383] = 25'b1101011110011111100011110;
      twice_table[384] = 25'b1101011110001000110111100;
      twice_table[385] = 25'b1101011101110010001100010;
      twice_table[386] = 25'b1101011101011011100010100;
      twice_table[387] = 25'b1101011101000100111001110;
      twice_table[388] = 25'b1101011100101110010010000;
      twice_table[389] = 25'b1101011100010111101011110;
      twice_table[390] = 25'b1101011100000001000110100;
      twice_table[391] = 25'b1101011011101010100010100;
      twice_table[392] = 25'b1101011011010011111111110;
      twice_table[393] = 25'b1101011010111101011110000;
      twice_table[394] = 25'b1101011010100110111101110;
      twice_table[395] = 25'b1101011010010000011110100;
      twice_table[396] = 25'b1101011001111010000000010;
      twice_table[397] = 25'b1101011001100011100011010;
      twice_table[398] = 25'b1101011001001101000111110;
      twice_table[399] = 25'b1101011000110110101101000;
      twice_table[400] = 25'b1101011000100000010011110;
      twice_table[401] = 25'b1101011000001001111011100;
      twice_table[402] = 25'b1101010111110011100100010;
      twice_table[403] = 25'b1101010111011101001110100;
      twice_table[404] = 25'b1101010111000110111001110;
      twice_table[405] = 25'b1101010110110000100110010;
      twice_table[406] = 25'b1101010110011010010011110;
      twice_table[407] = 25'b1101010110000100000010100;
      twice_table[408] = 25'b1101010101101101110010100;
      twice_table[409] = 25'b1101010101010111100011100;
      twice_table[410] = 25'b1101010101000001010101110;
      twice_table[411] = 25'b1101010100101011001001010;
      twice_table[412] = 25'b1101010100010100111101110;
      twice_table[413] = 25'b1101010011111110110011100;
      twice_table[414] = 25'b1101010011101000101010010;
      twice_table[415] = 25'b1101010011010010100010010;
      twice_table[416] = 25'b1101010010111100011011100;
      twice_table[417] = 25'b1101010010100110010101110;
      twice_table[418] = 25'b1101010010010000010001010;
      twice_table[419] = 25'b1101010001111010001101110;
      twice_table[420] = 25'b1101010001100100001011100;
      twice_table[421] = 25'b1101010001001110001010100;
      twice_table[422] = 25'b1101010000111000001010100;
      twice_table[423] = 25'b1101010000100010001011110;
      twice_table[424] = 25'b1101010000001100001110000;
      twice_table[425] = 25'b1101001111110110010001010;
      twice_table[426] = 25'b1101001111100000010110000;
      twice_table[427] = 25'b1101001111001010011011110;
      twice_table[428] = 25'b1101001110110100100010100;
      twice_table[429] = 25'b1101001110011110101010100;
      twice_table[430] = 25'b1101001110001000110011100;
      twice_table[431] = 25'b1101001101110010111101110;
      twice_table[432] = 25'b1101001101011101001001000;
      twice_table[433] = 25'b1101001101000111010101100;
      twice_table[434] = 25'b1101001100110001100011010;
      twice_table[435] = 25'b1101001100011011110010000;
      twice_table[436] = 25'b1101001100000110000001110;
      twice_table[437] = 25'b1101001011110000010010110;
      twice_table[438] = 25'b1101001011011010100100110;
      twice_table[439] = 25'b1101001011000100111000000;
      twice_table[440] = 25'b1101001010101111001100010;
      twice_table[441] = 25'b1101001010011001100001110;
      twice_table[442] = 25'b1101001010000011111000010;
      twice_table[443] = 25'b1101001001101110010000000;
      twice_table[444] = 25'b1101001001011000101000110;
      twice_table[445] = 25'b1101001001000011000010110;
      twice_table[446] = 25'b1101001000101101011101110;
      twice_table[447] = 25'b1101001000010111111001110;
      twice_table[448] = 25'b1101001000000010010111000;
      twice_table[449] = 25'b1101000111101100110101010;
      twice_table[450] = 25'b1101000111010111010100110;
      twice_table[451] = 25'b1101000111000001110101010;
      twice_table[452] = 25'b1101000110101100010110110;
      twice_table[453] = 25'b1101000110010110111001100;
      twice_table[454] = 25'b1101000110000001011101010;
      twice_table[455] = 25'b1101000101101100000010010;
      twice_table[456] = 25'b1101000101010110101000010;
      twice_table[457] = 25'b1101000101000001001111010;
      twice_table[458] = 25'b1101000100101011110111100;
      twice_table[459] = 25'b1101000100010110100000110;
      twice_table[460] = 25'b1101000100000001001011000;
      twice_table[461] = 25'b1101000011101011110110100;
      twice_table[462] = 25'b1101000011010110100011000;
      twice_table[463] = 25'b1101000011000001010000110;
      twice_table[464] = 25'b1101000010101011111111100;
      twice_table[465] = 25'b1101000010010110101111010;
      twice_table[466] = 25'b1101000010000001100000000;
      twice_table[467] = 25'b1101000001101100010010000;
      twice_table[468] = 25'b1101000001010111000101000;
      twice_table[469] = 25'b1101000001000001111001010;
      twice_table[470] = 25'b1101000000101100101110100;
      twice_table[471] = 25'b1101000000010111100100110;
      twice_table[472] = 25'b1101000000000010011100000;
      twice_table[473] = 25'b1100111111101101010100100;
      twice_table[474] = 25'b1100111111011000001110000;
      twice_table[475] = 25'b1100111111000011001000100;
      twice_table[476] = 25'b1100111110101110000100000;
      twice_table[477] = 25'b1100111110011001000000110;
      twice_table[478] = 25'b1100111110000011111110100;
      twice_table[479] = 25'b1100111101101110111101010;
      twice_table[480] = 25'b1100111101011001111101010;
      twice_table[481] = 25'b1100111101000100111110010;
      twice_table[482] = 25'b1100111100110000000000010;
      twice_table[483] = 25'b1100111100011011000011010;
      twice_table[484] = 25'b1100111100000110000111100;
      twice_table[485] = 25'b1100111011110001001100100;
      twice_table[486] = 25'b1100111011011100010010110;
      twice_table[487] = 25'b1100111011000111011010010;
      twice_table[488] = 25'b1100111010110010100010100;
      twice_table[489] = 25'b1100111010011101101100000;
      twice_table[490] = 25'b1100111010001000110110010;
      twice_table[491] = 25'b1100111001110100000001110;
      twice_table[492] = 25'b1100111001011111001110100;
      twice_table[493] = 25'b1100111001001010011100000;
      twice_table[494] = 25'b1100111000110101101010110;
      twice_table[495] = 25'b1100111000100000111010100;
      twice_table[496] = 25'b1100111000001100001011000;
      twice_table[497] = 25'b1100110111110111011101000;
      twice_table[498] = 25'b1100110111100010101111110;
      twice_table[499] = 25'b1100110111001110000011100;
      twice_table[500] = 25'b1100110110111001011000100;
      twice_table[501] = 25'b1100110110100100101110100;
      twice_table[502] = 25'b1100110110010000000101100;
      twice_table[503] = 25'b1100110101111011011101100;
      twice_table[504] = 25'b1100110101100110110110100;
      twice_table[505] = 25'b1100110101010010010000100;
      twice_table[506] = 25'b1100110100111101101011110;
      twice_table[507] = 25'b1100110100101001000111110;
      twice_table[508] = 25'b1100110100010100100101000;
      twice_table[509] = 25'b1100110100000000000011010;
      twice_table[510] = 25'b1100110011101011100010100;
      twice_table[511] = 25'b1100110011010111000010110;
      twice_table[512] = 25'b1100110011000010100100000;
      twice_table[513] = 25'b1100110010101110000110010;
      twice_table[514] = 25'b1100110010011001101001100;
      twice_table[515] = 25'b1100110010000101001110000;
      twice_table[516] = 25'b1100110001110000110011010;
      twice_table[517] = 25'b1100110001011100011001110;
      twice_table[518] = 25'b1100110001001000000001000;
      twice_table[519] = 25'b1100110000110011101001100;
      twice_table[520] = 25'b1100110000011111010011000;
      twice_table[521] = 25'b1100110000001010111101100;
      twice_table[522] = 25'b1100101111110110101000110;
      twice_table[523] = 25'b1100101111100010010101010;
      twice_table[524] = 25'b1100101111001110000010110;
      twice_table[525] = 25'b1100101110111001110001010;
      twice_table[526] = 25'b1100101110100101100000110;
      twice_table[527] = 25'b1100101110010001010001010;
      twice_table[528] = 25'b1100101101111101000010110;
      twice_table[529] = 25'b1100101101101000110101010;
      twice_table[530] = 25'b1100101101010100101000110;
      twice_table[531] = 25'b1100101101000000011101100;
      twice_table[532] = 25'b1100101100101100010011000;
      twice_table[533] = 25'b1100101100011000001001100;
      twice_table[534] = 25'b1100101100000100000001000;
      twice_table[535] = 25'b1100101011101111111001100;
      twice_table[536] = 25'b1100101011011011110011000;
      twice_table[537] = 25'b1100101011000111101101100;
      twice_table[538] = 25'b1100101010110011101001000;
      twice_table[539] = 25'b1100101010011111100101100;
      twice_table[540] = 25'b1100101010001011100011000;
      twice_table[541] = 25'b1100101001110111100001100;
      twice_table[542] = 25'b1100101001100011100001000;
      twice_table[543] = 25'b1100101001001111100001100;
      twice_table[544] = 25'b1100101000111011100010110;
      twice_table[545] = 25'b1100101000100111100101010;
      twice_table[546] = 25'b1100101000010011101000110;
      twice_table[547] = 25'b1100100111111111101101000;
      twice_table[548] = 25'b1100100111101011110010100;
      twice_table[549] = 25'b1100100111010111111000110;
      twice_table[550] = 25'b1100100111000100000000010;
      twice_table[551] = 25'b1100100110110000001000100;
      twice_table[552] = 25'b1100100110011100010001110;
      twice_table[553] = 25'b1100100110001000011100000;
      twice_table[554] = 25'b1100100101110100100111010;
      twice_table[555] = 25'b1100100101100000110011100;
      twice_table[556] = 25'b1100100101001101000000110;
      twice_table[557] = 25'b1100100100111001001111000;
      twice_table[558] = 25'b1100100100100101011110000;
      twice_table[559] = 25'b1100100100010001101110010;
      twice_table[560] = 25'b1100100011111101111111010;
      twice_table[561] = 25'b1100100011101010010001010;
      twice_table[562] = 25'b1100100011010110100100010;
      twice_table[563] = 25'b1100100011000010111000010;
      twice_table[564] = 25'b1100100010101111001101010;
      twice_table[565] = 25'b1100100010011011100011010;
      twice_table[566] = 25'b1100100010000111111010000;
      twice_table[567] = 25'b1100100001110100010001110;
      twice_table[568] = 25'b1100100001100000101010110;
      twice_table[569] = 25'b1100100001001101000100100;
      twice_table[570] = 25'b1100100000111001011111010;
      twice_table[571] = 25'b1100100000100101111010110;
      twice_table[572] = 25'b1100100000010010010111100;
      twice_table[573] = 25'b1100011111111110110101000;
      twice_table[574] = 25'b1100011111101011010011100;
      twice_table[575] = 25'b1100011111010111110011000;
      twice_table[576] = 25'b1100011111000100010011100;
      twice_table[577] = 25'b1100011110110000110100110;
      twice_table[578] = 25'b1100011110011101010111010;
      twice_table[579] = 25'b1100011110001001111010100;
      twice_table[580] = 25'b1100011101110110011110110;
      twice_table[581] = 25'b1100011101100011000100000;
      twice_table[582] = 25'b1100011101001111101010000;
      twice_table[583] = 25'b1100011100111100010001000;
      twice_table[584] = 25'b1100011100101000111001000;
      twice_table[585] = 25'b1100011100010101100010000;
      twice_table[586] = 25'b1100011100000010001100000;
      twice_table[587] = 25'b1100011011101110110110110;
      twice_table[588] = 25'b1100011011011011100010100;
      twice_table[589] = 25'b1100011011001000001111010;
      twice_table[590] = 25'b1100011010110100111101000;
      twice_table[591] = 25'b1100011010100001101011100;
      twice_table[592] = 25'b1100011010001110011011000;
      twice_table[593] = 25'b1100011001111011001011100;
      twice_table[594] = 25'b1100011001100111111100110;
      twice_table[595] = 25'b1100011001010100101111000;
      twice_table[596] = 25'b1100011001000001100010010;
      twice_table[597] = 25'b1100011000101110010110100;
      twice_table[598] = 25'b1100011000011011001011100;
      twice_table[599] = 25'b1100011000001000000001110;
      twice_table[600] = 25'b1100010111110100111000100;
      twice_table[601] = 25'b1100010111100001110000100;
      twice_table[602] = 25'b1100010111001110101001010;
      twice_table[603] = 25'b1100010110111011100011000;
      twice_table[604] = 25'b1100010110101000011101110;
      twice_table[605] = 25'b1100010110010101011001010;
      twice_table[606] = 25'b1100010110000010010101110;
      twice_table[607] = 25'b1100010101101111010011000;
      twice_table[608] = 25'b1100010101011100010001100;
      twice_table[609] = 25'b1100010101001001010000110;
      twice_table[610] = 25'b1100010100110110010000110;
      twice_table[611] = 25'b1100010100100011010001110;
      twice_table[612] = 25'b1100010100010000010011110;
      twice_table[613] = 25'b1100010011111101010110110;
      twice_table[614] = 25'b1100010011101010011010100;
      twice_table[615] = 25'b1100010011010111011111010;
      twice_table[616] = 25'b1100010011000100100100110;
      twice_table[617] = 25'b1100010010110001101011010;
      twice_table[618] = 25'b1100010010011110110010110;
      twice_table[619] = 25'b1100010010001011111011010;
      twice_table[620] = 25'b1100010001111001000100100;
      twice_table[621] = 25'b1100010001100110001110100;
      twice_table[622] = 25'b1100010001010011011001100;
      twice_table[623] = 25'b1100010001000000100101100;
      twice_table[624] = 25'b1100010000101101110010100;
      twice_table[625] = 25'b1100010000011011000000010;
      twice_table[626] = 25'b1100010000001000001110110;
      twice_table[627] = 25'b1100001111110101011110100;
      twice_table[628] = 25'b1100001111100010101110110;
      twice_table[629] = 25'b1100001111010000000000010;
      twice_table[630] = 25'b1100001110111101010010100;
      twice_table[631] = 25'b1100001110101010100101100;
      twice_table[632] = 25'b1100001110010111111001100;
      twice_table[633] = 25'b1100001110000101001110100;
      twice_table[634] = 25'b1100001101110010100100010;
      twice_table[635] = 25'b1100001101011111111011000;
      twice_table[636] = 25'b1100001101001101010010110;
      twice_table[637] = 25'b1100001100111010101011000;
      twice_table[638] = 25'b1100001100101000000100100;
      twice_table[639] = 25'b1100001100010101011110110;
      twice_table[640] = 25'b1100001100000010111001110;
      twice_table[641] = 25'b1100001011110000010110000;
      twice_table[642] = 25'b1100001011011101110010110;
      twice_table[643] = 25'b1100001011001011010000100;
      twice_table[644] = 25'b1100001010111000101111010;
      twice_table[645] = 25'b1100001010100110001110110;
      twice_table[646] = 25'b1100001010010011101111010;
      twice_table[647] = 25'b1100001010000001010000100;
      twice_table[648] = 25'b1100001001101110110010110;
      twice_table[649] = 25'b1100001001011100010101110;
      twice_table[650] = 25'b1100001001001001111001110;
      twice_table[651] = 25'b1100001000110111011110100;
      twice_table[652] = 25'b1100001000100101000100010;
      twice_table[653] = 25'b1100001000010010101010110;
      twice_table[654] = 25'b1100001000000000010010010;
      twice_table[655] = 25'b1100000111101101111010100;
      twice_table[656] = 25'b1100000111011011100011110;
      twice_table[657] = 25'b1100000111001001001101110;
      twice_table[658] = 25'b1100000110110110111000100;
      twice_table[659] = 25'b1100000110100100100100010;
      twice_table[660] = 25'b1100000110010010010001000;
      twice_table[661] = 25'b1100000101111111111110100;
      twice_table[662] = 25'b1100000101101101101100110;
      twice_table[663] = 25'b1100000101011011011100000;
      twice_table[664] = 25'b1100000101001001001100010;
      twice_table[665] = 25'b1100000100110110111101000;
      twice_table[666] = 25'b1100000100100100101111000;
      twice_table[667] = 25'b1100000100010010100001100;
      twice_table[668] = 25'b1100000100000000010101000;
      twice_table[669] = 25'b1100000011101110001001100;
      twice_table[670] = 25'b1100000011011011111110110;
      twice_table[671] = 25'b1100000011001001110100110;
      twice_table[672] = 25'b1100000010110111101011110;
      twice_table[673] = 25'b1100000010100101100011100;
      twice_table[674] = 25'b1100000010010011011100010;
      twice_table[675] = 25'b1100000010000001010101110;
      twice_table[676] = 25'b1100000001101111010000000;
      twice_table[677] = 25'b1100000001011101001011010;
      twice_table[678] = 25'b1100000001001011000111010;
      twice_table[679] = 25'b1100000000111001000100010;
      twice_table[680] = 25'b1100000000100111000010000;
      twice_table[681] = 25'b1100000000010101000000100;
      twice_table[682] = 25'b1100000000000011000000000;
      twice_table[683] = 25'b1011111111110001000000010;
      twice_table[684] = 25'b1011111111011111000001100;
      twice_table[685] = 25'b1011111111001101000011100;
      twice_table[686] = 25'b1011111110111011000110010;
      twice_table[687] = 25'b1011111110101001001001110;
      twice_table[688] = 25'b1011111110010111001110010;
      twice_table[689] = 25'b1011111110000101010011110;
      twice_table[690] = 25'b1011111101110011011001110;
      twice_table[691] = 25'b1011111101100001100000110;
      twice_table[692] = 25'b1011111101001111101000110;
      twice_table[693] = 25'b1011111100111101110001010;
      twice_table[694] = 25'b1011111100101011111010110;
      twice_table[695] = 25'b1011111100011010000101010;
      twice_table[696] = 25'b1011111100001000010000010;
      twice_table[697] = 25'b1011111011110110011100010;
      twice_table[698] = 25'b1011111011100100101001010;
      twice_table[699] = 25'b1011111011010010110110110;
      twice_table[700] = 25'b1011111011000001000101010;
      twice_table[701] = 25'b1011111010101111010100100;
      twice_table[702] = 25'b1011111010011101100100110;
      twice_table[703] = 25'b1011111010001011110101110;
      twice_table[704] = 25'b1011111001111010000111100;
      twice_table[705] = 25'b1011111001101000011010010;
      twice_table[706] = 25'b1011111001010110101101100;
      twice_table[707] = 25'b1011111001000101000001110;
      twice_table[708] = 25'b1011111000110011010111000;
      twice_table[709] = 25'b1011111000100001101100110;
      twice_table[710] = 25'b1011111000010000000011100;
      twice_table[711] = 25'b1011110111111110011011000;
      twice_table[712] = 25'b1011110111101100110011100;
      twice_table[713] = 25'b1011110111011011001100100;
      twice_table[714] = 25'b1011110111001001100110100;
      twice_table[715] = 25'b1011110110111000000001100;
      twice_table[716] = 25'b1011110110100110011101000;
      twice_table[717] = 25'b1011110110010100111001100;
      twice_table[718] = 25'b1011110110000011010110110;
      twice_table[719] = 25'b1011110101110001110100110;
      twice_table[720] = 25'b1011110101100000010011100;
      twice_table[721] = 25'b1011110101001110110011010;
      twice_table[722] = 25'b1011110100111101010011110;
      twice_table[723] = 25'b1011110100101011110101000;
      twice_table[724] = 25'b1011110100011010010111010;
      twice_table[725] = 25'b1011110100001000111010000;
      twice_table[726] = 25'b1011110011110111011101110;
      twice_table[727] = 25'b1011110011100110000010010;
      twice_table[728] = 25'b1011110011010100100111100;
      twice_table[729] = 25'b1011110011000011001101110;
      twice_table[730] = 25'b1011110010110001110100110;
      twice_table[731] = 25'b1011110010100000011100010;
      twice_table[732] = 25'b1011110010001111000101000;
      twice_table[733] = 25'b1011110001111101101110010;
      twice_table[734] = 25'b1011110001101100011000010;
      twice_table[735] = 25'b1011110001011011000011010;
      twice_table[736] = 25'b1011110001001001101111000;
      twice_table[737] = 25'b1011110000111000011011100;
      twice_table[738] = 25'b1011110000100111001000110;
      twice_table[739] = 25'b1011110000010101110111000;
      twice_table[740] = 25'b1011110000000100100101110;
      twice_table[741] = 25'b1011101111110011010101100;
      twice_table[742] = 25'b1011101111100010000110000;
      twice_table[743] = 25'b1011101111010000110111010;
      twice_table[744] = 25'b1011101110111111101001010;
      twice_table[745] = 25'b1011101110101110011100000;
      twice_table[746] = 25'b1011101110011101001111110;
      twice_table[747] = 25'b1011101110001100000100010;
      twice_table[748] = 25'b1011101101111010111001010;
      twice_table[749] = 25'b1011101101101001101111010;
      twice_table[750] = 25'b1011101101011000100110010;
      twice_table[751] = 25'b1011101101000111011101110;
      twice_table[752] = 25'b1011101100110110010110000;
      twice_table[753] = 25'b1011101100100101001111010;
      twice_table[754] = 25'b1011101100010100001001000;
      twice_table[755] = 25'b1011101100000011000011110;
      twice_table[756] = 25'b1011101011110001111111010;
      twice_table[757] = 25'b1011101011100000111011100;
      twice_table[758] = 25'b1011101011001111111000100;
      twice_table[759] = 25'b1011101010111110110110010;
      twice_table[760] = 25'b1011101010101101110101000;
      twice_table[761] = 25'b1011101010011100110100010;
      twice_table[762] = 25'b1011101010001011110100100;
      twice_table[763] = 25'b1011101001111010110101010;
      twice_table[764] = 25'b1011101001101001110111000;
      twice_table[765] = 25'b1011101001011000111001100;
      twice_table[766] = 25'b1011101001000111111100110;
      twice_table[767] = 25'b1011101000110111000000110;
      twice_table[768] = 25'b1011101000100110000101100;
      twice_table[769] = 25'b1011101000010101001011000;
      twice_table[770] = 25'b1011101000000100010001010;
      twice_table[771] = 25'b1011100111110011011000010;
      twice_table[772] = 25'b1011100111100010100000000;
      twice_table[773] = 25'b1011100111010001101000110;
      twice_table[774] = 25'b1011100111000000110010000;
      twice_table[775] = 25'b1011100110101111111100010;
      twice_table[776] = 25'b1011100110011111000111000;
      twice_table[777] = 25'b1011100110001110010010110;
      twice_table[778] = 25'b1011100101111101011111010;
      twice_table[779] = 25'b1011100101101100101100010;
      twice_table[780] = 25'b1011100101011011111010010;
      twice_table[781] = 25'b1011100101001011001001000;
      twice_table[782] = 25'b1011100100111010011000100;
      twice_table[783] = 25'b1011100100101001101000100;
      twice_table[784] = 25'b1011100100011000111001100;
      twice_table[785] = 25'b1011100100001000001011010;
      twice_table[786] = 25'b1011100011110111011101110;
      twice_table[787] = 25'b1011100011100110110001000;
      twice_table[788] = 25'b1011100011010110000101000;
      twice_table[789] = 25'b1011100011000101011001110;
      twice_table[790] = 25'b1011100010110100101111010;
      twice_table[791] = 25'b1011100010100100000101100;
      twice_table[792] = 25'b1011100010010011011100100;
      twice_table[793] = 25'b1011100010000010110100010;
      twice_table[794] = 25'b1011100001110010001100110;
      twice_table[795] = 25'b1011100001100001100110000;
      twice_table[796] = 25'b1011100001010001000000000;
      twice_table[797] = 25'b1011100001000000011010110;
      twice_table[798] = 25'b1011100000101111110110000;
      twice_table[799] = 25'b1011100000011111010010010;
      twice_table[800] = 25'b1011100000001110101111010;
      twice_table[801] = 25'b1011011111111110001101000;
      twice_table[802] = 25'b1011011111101101101011100;
      twice_table[803] = 25'b1011011111011101001010110;
      twice_table[804] = 25'b1011011111001100101010100;
      twice_table[805] = 25'b1011011110111100001011010;
      twice_table[806] = 25'b1011011110101011101100110;
      twice_table[807] = 25'b1011011110011011001110110;
      twice_table[808] = 25'b1011011110001010110001110;
      twice_table[809] = 25'b1011011101111010010101010;
      twice_table[810] = 25'b1011011101101001111001110;
      twice_table[811] = 25'b1011011101011001011110110;
      twice_table[812] = 25'b1011011101001001000100110;
      twice_table[813] = 25'b1011011100111000101011010;
      twice_table[814] = 25'b1011011100101000010010100;
      twice_table[815] = 25'b1011011100010111111010100;
      twice_table[816] = 25'b1011011100000111100011010;
      twice_table[817] = 25'b1011011011110111001100110;
      twice_table[818] = 25'b1011011011100110110111000;
      twice_table[819] = 25'b1011011011010110100010000;
      twice_table[820] = 25'b1011011011000110001101110;
      twice_table[821] = 25'b1011011010110101111010000;
      twice_table[822] = 25'b1011011010100101100111010;
      twice_table[823] = 25'b1011011010010101010101000;
      twice_table[824] = 25'b1011011010000101000011110;
      twice_table[825] = 25'b1011011001110100110011000;
      twice_table[826] = 25'b1011011001100100100011000;
      twice_table[827] = 25'b1011011001010100010011110;
      twice_table[828] = 25'b1011011001000100000101010;
      twice_table[829] = 25'b1011011000110011110111100;
      twice_table[830] = 25'b1011011000100011101010100;
      twice_table[831] = 25'b1011011000010011011110000;
      twice_table[832] = 25'b1011011000000011010010100;
      twice_table[833] = 25'b1011010111110011000111100;
      twice_table[834] = 25'b1011010111100010111101010;
      twice_table[835] = 25'b1011010111010010110011110;
      twice_table[836] = 25'b1011010111000010101011000;
      twice_table[837] = 25'b1011010110110010100011000;
      twice_table[838] = 25'b1011010110100010011011110;
      twice_table[839] = 25'b1011010110010010010101000;
      twice_table[840] = 25'b1011010110000010001111010;
      twice_table[841] = 25'b1011010101110010001010000;
      twice_table[842] = 25'b1011010101100010000101100;
      twice_table[843] = 25'b1011010101010010000001110;
      twice_table[844] = 25'b1011010101000001111110110;
      twice_table[845] = 25'b1011010100110001111100100;
      twice_table[846] = 25'b1011010100100001111010110;
      twice_table[847] = 25'b1011010100010001111001110;
      twice_table[848] = 25'b1011010100000001111001100;
      twice_table[849] = 25'b1011010011110001111010000;
      twice_table[850] = 25'b1011010011100001111011010;
      twice_table[851] = 25'b1011010011010001111101010;
      twice_table[852] = 25'b1011010011000001111111110;
      twice_table[853] = 25'b1011010010110010000011000;
      twice_table[854] = 25'b1011010010100010000111000;
      twice_table[855] = 25'b1011010010010010001011110;
      twice_table[856] = 25'b1011010010000010010001010;
      twice_table[857] = 25'b1011010001110010010111010;
      twice_table[858] = 25'b1011010001100010011110010;
      twice_table[859] = 25'b1011010001010010100101110;
      twice_table[860] = 25'b1011010001000010101110000;
      twice_table[861] = 25'b1011010000110010110110110;
      twice_table[862] = 25'b1011010000100011000000100;
      twice_table[863] = 25'b1011010000010011001010110;
      twice_table[864] = 25'b1011010000000011010101110;
      twice_table[865] = 25'b1011001111110011100001100;
      twice_table[866] = 25'b1011001111100011101101110;
      twice_table[867] = 25'b1011001111010011111011000;
      twice_table[868] = 25'b1011001111000100001000110;
      twice_table[869] = 25'b1011001110110100010111010;
      twice_table[870] = 25'b1011001110100100100110100;
      twice_table[871] = 25'b1011001110010100110110010;
      twice_table[872] = 25'b1011001110000101000110110;
      twice_table[873] = 25'b1011001101110101011000000;
      twice_table[874] = 25'b1011001101100101101010000;
      twice_table[875] = 25'b1011001101010101111100100;
      twice_table[876] = 25'b1011001101000110001111110;
      twice_table[877] = 25'b1011001100110110100011110;
      twice_table[878] = 25'b1011001100100110111000100;
      twice_table[879] = 25'b1011001100010111001110000;
      twice_table[880] = 25'b1011001100000111100100000;
      twice_table[881] = 25'b1011001011110111111010110;
      twice_table[882] = 25'b1011001011101000010010000;
      twice_table[883] = 25'b1011001011011000101010010;
      twice_table[884] = 25'b1011001011001001000011000;
      twice_table[885] = 25'b1011001010111001011100100;
      twice_table[886] = 25'b1011001010101001110110100;
      twice_table[887] = 25'b1011001010011010010001100;
      twice_table[888] = 25'b1011001010001010101101000;
      twice_table[889] = 25'b1011001001111011001001000;
      twice_table[890] = 25'b1011001001101011100110000;
      twice_table[891] = 25'b1011001001011100000011100;
      twice_table[892] = 25'b1011001001001100100001110;
      twice_table[893] = 25'b1011001000111101000000100;
      twice_table[894] = 25'b1011001000101101100000000;
      twice_table[895] = 25'b1011001000011110000000010;
      twice_table[896] = 25'b1011001000001110100001010;
      twice_table[897] = 25'b1011000111111111000010110;
      twice_table[898] = 25'b1011000111101111100101000;
      twice_table[899] = 25'b1011000111100000001000000;
      twice_table[900] = 25'b1011000111010000101011100;
      twice_table[901] = 25'b1011000111000001001111110;
      twice_table[902] = 25'b1011000110110001110100110;
      twice_table[903] = 25'b1011000110100010011010100;
      twice_table[904] = 25'b1011000110010011000000110;
      twice_table[905] = 25'b1011000110000011100111100;
      twice_table[906] = 25'b1011000101110100001111010;
      twice_table[907] = 25'b1011000101100100110111100;
      twice_table[908] = 25'b1011000101010101100000100;
      twice_table[909] = 25'b1011000101000110001010000;
      twice_table[910] = 25'b1011000100110110110100010;
      twice_table[911] = 25'b1011000100100111011111010;
      twice_table[912] = 25'b1011000100011000001010110;
      twice_table[913] = 25'b1011000100001000110111000;
      twice_table[914] = 25'b1011000011111001100100000;
      twice_table[915] = 25'b1011000011101010010001100;
      twice_table[916] = 25'b1011000011011010111111110;
      twice_table[917] = 25'b1011000011001011101110110;
      twice_table[918] = 25'b1011000010111100011110010;
      twice_table[919] = 25'b1011000010101101001110100;
      twice_table[920] = 25'b1011000010011101111111010;
      twice_table[921] = 25'b1011000010001110110000110;
      twice_table[922] = 25'b1011000001111111100011000;
      twice_table[923] = 25'b1011000001110000010110000;
      twice_table[924] = 25'b1011000001100001001001100;
      twice_table[925] = 25'b1011000001010001111101100;
      twice_table[926] = 25'b1011000001000010110010010;
      twice_table[927] = 25'b1011000000110011100111110;
      twice_table[928] = 25'b1011000000100100011110000;
      twice_table[929] = 25'b1011000000010101010100110;
      twice_table[930] = 25'b1011000000000110001100000;
      twice_table[931] = 25'b1010111111110111000100000;
      twice_table[932] = 25'b1010111111100111111100110;
      twice_table[933] = 25'b1010111111011000110110010;
      twice_table[934] = 25'b1010111111001001110000010;
      twice_table[935] = 25'b1010111110111010101010110;
      twice_table[936] = 25'b1010111110101011100110010;
      twice_table[937] = 25'b1010111110011100100010000;
      twice_table[938] = 25'b1010111110001101011110110;
      twice_table[939] = 25'b1010111101111110011100000;
      twice_table[940] = 25'b1010111101101111011001110;
      twice_table[941] = 25'b1010111101100000011000010;
      twice_table[942] = 25'b1010111101010001010111100;
      twice_table[943] = 25'b1010111101000010010111010;
      twice_table[944] = 25'b1010111100110011010111110;
      twice_table[945] = 25'b1010111100100100011000110;
      twice_table[946] = 25'b1010111100010101011010100;
      twice_table[947] = 25'b1010111100000110011101000;
      twice_table[948] = 25'b1010111011110111100000000;
      twice_table[949] = 25'b1010111011101000100011100;
      twice_table[950] = 25'b1010111011011001101000000;
      twice_table[951] = 25'b1010111011001010101100110;
      twice_table[952] = 25'b1010111010111011110010100;
      twice_table[953] = 25'b1010111010101100111000100;
      twice_table[954] = 25'b1010111010011101111111100;
      twice_table[955] = 25'b1010111010001111000111000;
      twice_table[956] = 25'b1010111010000000001111000;
      twice_table[957] = 25'b1010111001110001010111110;
      twice_table[958] = 25'b1010111001100010100001000;
      twice_table[959] = 25'b1010111001010011101011000;
      twice_table[960] = 25'b1010111001000100110101110;
      twice_table[961] = 25'b1010111000110110000001000;
      twice_table[962] = 25'b1010111000100111001101000;
      twice_table[963] = 25'b1010111000011000011001100;
      twice_table[964] = 25'b1010111000001001100110100;
      twice_table[965] = 25'b1010110111111010110100010;
      twice_table[966] = 25'b1010110111101100000010110;
      twice_table[967] = 25'b1010110111011101010001110;
      twice_table[968] = 25'b1010110111001110100001100;
      twice_table[969] = 25'b1010110110111111110001110;
      twice_table[970] = 25'b1010110110110001000010110;
      twice_table[971] = 25'b1010110110100010010100010;
      twice_table[972] = 25'b1010110110010011100110010;
      twice_table[973] = 25'b1010110110000100111001010;
      twice_table[974] = 25'b1010110101110110001100100;
      twice_table[975] = 25'b1010110101100111100000100;
      twice_table[976] = 25'b1010110101011000110101010;
      twice_table[977] = 25'b1010110101001010001010100;
      twice_table[978] = 25'b1010110100111011100000100;
      twice_table[979] = 25'b1010110100101100110111000;
      twice_table[980] = 25'b1010110100011110001110000;
      twice_table[981] = 25'b1010110100001111100101110;
      twice_table[982] = 25'b1010110100000000111110010;
      twice_table[983] = 25'b1010110011110010010111010;
      twice_table[984] = 25'b1010110011100011110000110;
      twice_table[985] = 25'b1010110011010101001011000;
      twice_table[986] = 25'b1010110011000110100101110;
      twice_table[987] = 25'b1010110010111000000001010;
      twice_table[988] = 25'b1010110010101001011101010;
      twice_table[989] = 25'b1010110010011010111010000;
      twice_table[990] = 25'b1010110010001100010111010;
      twice_table[991] = 25'b1010110001111101110101010;
      twice_table[992] = 25'b1010110001101111010011110;
      twice_table[993] = 25'b1010110001100000110010110;
      twice_table[994] = 25'b1010110001010010010010100;
      twice_table[995] = 25'b1010110001000011110011000;
      twice_table[996] = 25'b1010110000110101010100000;
      twice_table[997] = 25'b1010110000100110110101100;
      twice_table[998] = 25'b1010110000011000010111100;
      twice_table[999] = 25'b1010110000001001111010100;
      twice_table[1000] = 25'b1010101111111011011101110;
      twice_table[1001] = 25'b1010101111101101000001110;
      twice_table[1002] = 25'b1010101111011110100110010;
      twice_table[1003] = 25'b1010101111010000001011100;
      twice_table[1004] = 25'b1010101111000001110001100;
      twice_table[1005] = 25'b1010101110110011010111110;
      twice_table[1006] = 25'b1010101110100100111110110;
      twice_table[1007] = 25'b1010101110010110100110100;
      twice_table[1008] = 25'b1010101110001000001110110;
      twice_table[1009] = 25'b1010101101111001110111100;
      twice_table[1010] = 25'b1010101101101011100001000;
      twice_table[1011] = 25'b1010101101011101001011000;
      twice_table[1012] = 25'b1010101101001110110101100;
      twice_table[1013] = 25'b1010101101000000100000110;
      twice_table[1014] = 25'b1010101100110010001100100;
      twice_table[1015] = 25'b1010101100100011111001000;
      twice_table[1016] = 25'b1010101100010101100110000;
      twice_table[1017] = 25'b1010101100000111010011110;
      twice_table[1018] = 25'b1010101011111001000001110;
      twice_table[1019] = 25'b1010101011101010110000110;
      twice_table[1020] = 25'b1010101011011100100000000;
      twice_table[1021] = 25'b1010101011001110010000000;
      twice_table[1022] = 25'b1010101011000000000000110;
      twice_table[1023] = 25'b1010101010110001110001110;
      twice_table[1024] = 25'b1010101010100011100011110;
      twice_table[1025] = 25'b1010101010010101010110000;
      twice_table[1026] = 25'b1010101010000111001001000;
      twice_table[1027] = 25'b1010101001111000111100100;
      twice_table[1028] = 25'b1010101001101010110000110;
      twice_table[1029] = 25'b1010101001011100100101100;
      twice_table[1030] = 25'b1010101001001110011010110;
      twice_table[1031] = 25'b1010101001000000010000110;
      twice_table[1032] = 25'b1010101000110010000111010;
      twice_table[1033] = 25'b1010101000100011111110010;
      twice_table[1034] = 25'b1010101000010101110110000;
      twice_table[1035] = 25'b1010101000000111101110010;
      twice_table[1036] = 25'b1010100111111001100111000;
      twice_table[1037] = 25'b1010100111101011100000100;
      twice_table[1038] = 25'b1010100111011101011010100;
      twice_table[1039] = 25'b1010100111001111010101000;
      twice_table[1040] = 25'b1010100111000001010000010;
      twice_table[1041] = 25'b1010100110110011001100000;
      twice_table[1042] = 25'b1010100110100101001000010;
      twice_table[1043] = 25'b1010100110010111000101010;
      twice_table[1044] = 25'b1010100110001001000010110;
      twice_table[1045] = 25'b1010100101111011000001000;
      twice_table[1046] = 25'b1010100101101100111111100;
      twice_table[1047] = 25'b1010100101011110111110110;
      twice_table[1048] = 25'b1010100101010000111110110;
      twice_table[1049] = 25'b1010100101000010111111000;
      twice_table[1050] = 25'b1010100100110101000000000;
      twice_table[1051] = 25'b1010100100100111000001110;
      twice_table[1052] = 25'b1010100100011001000011110;
      twice_table[1053] = 25'b1010100100001011000110100;
      twice_table[1054] = 25'b1010100011111101001001110;
      twice_table[1055] = 25'b1010100011101111001101110;
      twice_table[1056] = 25'b1010100011100001010010010;
      twice_table[1057] = 25'b1010100011010011010111010;
      twice_table[1058] = 25'b1010100011000101011100110;
      twice_table[1059] = 25'b1010100010110111100011000;
      twice_table[1060] = 25'b1010100010101001101001110;
      twice_table[1061] = 25'b1010100010011011110001000;
      twice_table[1062] = 25'b1010100010001101111000110;
      twice_table[1063] = 25'b1010100010000000000001010;
      twice_table[1064] = 25'b1010100001110010001010010;
      twice_table[1065] = 25'b1010100001100100010100000;
      twice_table[1066] = 25'b1010100001010110011110000;
      twice_table[1067] = 25'b1010100001001000101000110;
      twice_table[1068] = 25'b1010100000111010110100010;
      twice_table[1069] = 25'b1010100000101101000000000;
      twice_table[1070] = 25'b1010100000011111001100100;
      twice_table[1071] = 25'b1010100000010001011001100;
      twice_table[1072] = 25'b1010100000000011100111000;
      twice_table[1073] = 25'b1010011111110101110101010;
      twice_table[1074] = 25'b1010011111101000000011110;
      twice_table[1075] = 25'b1010011111011010010011000;
      twice_table[1076] = 25'b1010011111001100100011000;
      twice_table[1077] = 25'b1010011110111110110011010;
      twice_table[1078] = 25'b1010011110110001000100010;
      twice_table[1079] = 25'b1010011110100011010101110;
      twice_table[1080] = 25'b1010011110010101101000000;
      twice_table[1081] = 25'b1010011110000111111010100;
      twice_table[1082] = 25'b1010011101111010001101110;
      twice_table[1083] = 25'b1010011101101100100001100;
      twice_table[1084] = 25'b1010011101011110110101110;
      twice_table[1085] = 25'b1010011101010001001010110;
      twice_table[1086] = 25'b1010011101000011100000000;
      twice_table[1087] = 25'b1010011100110101110110000;
      twice_table[1088] = 25'b1010011100101000001100110;
      twice_table[1089] = 25'b1010011100011010100011110;
      twice_table[1090] = 25'b1010011100001100111011100;
      twice_table[1091] = 25'b1010011011111111010011110;
      twice_table[1092] = 25'b1010011011110001101100100;
      twice_table[1093] = 25'b1010011011100100000101110;
      twice_table[1094] = 25'b1010011011010110011111110;
      twice_table[1095] = 25'b1010011011001000111010000;
      twice_table[1096] = 25'b1010011010111011010101000;
      twice_table[1097] = 25'b1010011010101101110000100;
      twice_table[1098] = 25'b1010011010100000001100110;
      twice_table[1099] = 25'b1010011010010010101001010;
      twice_table[1100] = 25'b1010011010000101000110100;
      twice_table[1101] = 25'b1010011001110111100100010;
      twice_table[1102] = 25'b1010011001101010000010100;
      twice_table[1103] = 25'b1010011001011100100001100;
      twice_table[1104] = 25'b1010011001001111000000110;
      twice_table[1105] = 25'b1010011001000001100000110;
      twice_table[1106] = 25'b1010011000110100000001010;
      twice_table[1107] = 25'b1010011000100110100010010;
      twice_table[1108] = 25'b1010011000011001000100000;
      twice_table[1109] = 25'b1010011000001011100110000;
      twice_table[1110] = 25'b1010010111111110001000110;
      twice_table[1111] = 25'b1010010111110000101100000;
      twice_table[1112] = 25'b1010010111100011001111110;
      twice_table[1113] = 25'b1010010111010101110100000;
      twice_table[1114] = 25'b1010010111001000011000110;
      twice_table[1115] = 25'b1010010110111010111110010;
      twice_table[1116] = 25'b1010010110101101100100010;
      twice_table[1117] = 25'b1010010110100000001010110;
      twice_table[1118] = 25'b1010010110010010110001110;
      twice_table[1119] = 25'b1010010110000101011001010;
      twice_table[1120] = 25'b1010010101111000000001010;
      twice_table[1121] = 25'b1010010101101010101010000;
      twice_table[1122] = 25'b1010010101011101010011010;
      twice_table[1123] = 25'b1010010101001111111101000;
      twice_table[1124] = 25'b1010010101000010100111010;
      twice_table[1125] = 25'b1010010100110101010010000;
      twice_table[1126] = 25'b1010010100100111111101010;
      twice_table[1127] = 25'b1010010100011010101001010;
      twice_table[1128] = 25'b1010010100001101010101110;
      twice_table[1129] = 25'b1010010100000000000010100;
      twice_table[1130] = 25'b1010010011110010110000000;
      twice_table[1131] = 25'b1010010011100101011110000;
      twice_table[1132] = 25'b1010010011011000001100110;
      twice_table[1133] = 25'b1010010011001010111011110;
      twice_table[1134] = 25'b1010010010111101101011010;
      twice_table[1135] = 25'b1010010010110000011011100;
      twice_table[1136] = 25'b1010010010100011001100010;
      twice_table[1137] = 25'b1010010010010101111101100;
      twice_table[1138] = 25'b1010010010001000101111010;
      twice_table[1139] = 25'b1010010001111011100001100;
      twice_table[1140] = 25'b1010010001101110010100010;
      twice_table[1141] = 25'b1010010001100001000111100;
      twice_table[1142] = 25'b1010010001010011111011100;
      twice_table[1143] = 25'b1010010001000110101111110;
      twice_table[1144] = 25'b1010010000111001100100110;
      twice_table[1145] = 25'b1010010000101100011010010;
      twice_table[1146] = 25'b1010010000011111010000010;
      twice_table[1147] = 25'b1010010000010010000110110;
      twice_table[1148] = 25'b1010010000000100111101110;
      twice_table[1149] = 25'b1010001111110111110101010;
      twice_table[1150] = 25'b1010001111101010101101100;
      twice_table[1151] = 25'b1010001111011101100110000;
      twice_table[1152] = 25'b1010001111010000011111010;
      twice_table[1153] = 25'b1010001111000011011000110;
      twice_table[1154] = 25'b1010001110110110010011000;
      twice_table[1155] = 25'b1010001110101001001101110;
      twice_table[1156] = 25'b1010001110011100001001000;
      twice_table[1157] = 25'b1010001110001111000100110;
      twice_table[1158] = 25'b1010001110000010000001000;
      twice_table[1159] = 25'b1010001101110100111101110;
      twice_table[1160] = 25'b1010001101100111111011010;
      twice_table[1161] = 25'b1010001101011010111001000;
      twice_table[1162] = 25'b1010001101001101110111010;
      twice_table[1163] = 25'b1010001101000000110110010;
      twice_table[1164] = 25'b1010001100110011110101100;
      twice_table[1165] = 25'b1010001100100110110101100;
      twice_table[1166] = 25'b1010001100011001110110000;
      twice_table[1167] = 25'b1010001100001100110111000;
      twice_table[1168] = 25'b1010001011111111111000010;
      twice_table[1169] = 25'b1010001011110010111010010;
      twice_table[1170] = 25'b1010001011100101111100110;
      twice_table[1171] = 25'b1010001011011000111111110;
      twice_table[1172] = 25'b1010001011001100000011100;
      twice_table[1173] = 25'b1010001010111111000111100;
      twice_table[1174] = 25'b1010001010110010001100000;
      twice_table[1175] = 25'b1010001010100101010001000;
      twice_table[1176] = 25'b1010001010011000010110110;
      twice_table[1177] = 25'b1010001010001011011100110;
      twice_table[1178] = 25'b1010001001111110100011010;
      twice_table[1179] = 25'b1010001001110001101010100;
      twice_table[1180] = 25'b1010001001100100110010000;
      twice_table[1181] = 25'b1010001001010111111010010;
      twice_table[1182] = 25'b1010001001001011000010110;
      twice_table[1183] = 25'b1010001000111110001100000;
      twice_table[1184] = 25'b1010001000110001010101110;
      twice_table[1185] = 25'b1010001000100100011111110;
      twice_table[1186] = 25'b1010001000010111101010100;
      twice_table[1187] = 25'b1010001000001010110101110;
      twice_table[1188] = 25'b1010000111111110000001100;
      twice_table[1189] = 25'b1010000111110001001101110;
      twice_table[1190] = 25'b1010000111100100011010010;
      twice_table[1191] = 25'b1010000111010111100111100;
      twice_table[1192] = 25'b1010000111001010110101010;
      twice_table[1193] = 25'b1010000110111110000011100;
      twice_table[1194] = 25'b1010000110110001010010010;
      twice_table[1195] = 25'b1010000110100100100001100;
      twice_table[1196] = 25'b1010000110010111110001010;
      twice_table[1197] = 25'b1010000110001011000001100;
      twice_table[1198] = 25'b1010000101111110010010010;
      twice_table[1199] = 25'b1010000101110001100011100;
      twice_table[1200] = 25'b1010000101100100110101010;
      twice_table[1201] = 25'b1010000101011000000111100;
      twice_table[1202] = 25'b1010000101001011011010010;
      twice_table[1203] = 25'b1010000100111110101101100;
      twice_table[1204] = 25'b1010000100110010000001010;
      twice_table[1205] = 25'b1010000100100101010101100;
      twice_table[1206] = 25'b1010000100011000101010010;
      twice_table[1207] = 25'b1010000100001011111111100;
      twice_table[1208] = 25'b1010000011111111010101010;
      twice_table[1209] = 25'b1010000011110010101011100;
      twice_table[1210] = 25'b1010000011100110000010010;
      twice_table[1211] = 25'b1010000011011001011001100;
      twice_table[1212] = 25'b1010000011001100110001010;
      twice_table[1213] = 25'b1010000011000000001001100;
      twice_table[1214] = 25'b1010000010110011100010010;
      twice_table[1215] = 25'b1010000010100110111011010;
      twice_table[1216] = 25'b1010000010011010010101000;
      twice_table[1217] = 25'b1010000010001101101111010;
      twice_table[1218] = 25'b1010000010000001001010000;
      twice_table[1219] = 25'b1010000001110100100101010;
      twice_table[1220] = 25'b1010000001101000000000110;
      twice_table[1221] = 25'b1010000001011011011101000;
      twice_table[1222] = 25'b1010000001001110111001110;
      twice_table[1223] = 25'b1010000001000010010110110;
      twice_table[1224] = 25'b1010000000110101110100100;
      twice_table[1225] = 25'b1010000000101001010010110;
      twice_table[1226] = 25'b1010000000011100110001010;
      twice_table[1227] = 25'b1010000000010000010000100;
      twice_table[1228] = 25'b1010000000000011110000000;
      twice_table[1229] = 25'b1001111111110111010000000;
      twice_table[1230] = 25'b1001111111101010110000110;
      twice_table[1231] = 25'b1001111111011110010001110;
      twice_table[1232] = 25'b1001111111010001110011010;
      twice_table[1233] = 25'b1001111111000101010101100;
      twice_table[1234] = 25'b1001111110111000111000000;
      twice_table[1235] = 25'b1001111110101100011011000;
      twice_table[1236] = 25'b1001111110011111111110100;
      twice_table[1237] = 25'b1001111110010011100010100;
      twice_table[1238] = 25'b1001111110000111000111000;
      twice_table[1239] = 25'b1001111101111010101011110;
      twice_table[1240] = 25'b1001111101101110010001010;
      twice_table[1241] = 25'b1001111101100001110111010;
      twice_table[1242] = 25'b1001111101010101011101110;
      twice_table[1243] = 25'b1001111101001001000100100;
      twice_table[1244] = 25'b1001111100111100101100000;
      twice_table[1245] = 25'b1001111100110000010011110;
      twice_table[1246] = 25'b1001111100100011111100000;
      twice_table[1247] = 25'b1001111100010111100101000;
      twice_table[1248] = 25'b1001111100001011001110010;
      twice_table[1249] = 25'b1001111011111110111000000;
      twice_table[1250] = 25'b1001111011110010100010010;
      twice_table[1251] = 25'b1001111011100110001101000;
      twice_table[1252] = 25'b1001111011011001111000010;
      twice_table[1253] = 25'b1001111011001101100011110;
      twice_table[1254] = 25'b1001111011000001010000000;
      twice_table[1255] = 25'b1001111010110100111100110;
      twice_table[1256] = 25'b1001111010101000101001110;
      twice_table[1257] = 25'b1001111010011100010111010;
      twice_table[1258] = 25'b1001111010010000000101100;
      twice_table[1259] = 25'b1001111010000011110100000;
      twice_table[1260] = 25'b1001111001110111100011000;
      twice_table[1261] = 25'b1001111001101011010010100;
      twice_table[1262] = 25'b1001111001011111000010100;
      twice_table[1263] = 25'b1001111001010010110011000;
      twice_table[1264] = 25'b1001111001000110100011110;
      twice_table[1265] = 25'b1001111000111010010101010;
      twice_table[1266] = 25'b1001111000101110000111000;
      twice_table[1267] = 25'b1001111000100001111001100;
      twice_table[1268] = 25'b1001111000010101101100010;
      twice_table[1269] = 25'b1001111000001001011111100;
      twice_table[1270] = 25'b1001110111111101010011010;
      twice_table[1271] = 25'b1001110111110001000111100;
      twice_table[1272] = 25'b1001110111100100111100000;
      twice_table[1273] = 25'b1001110111011000110001010;
      twice_table[1274] = 25'b1001110111001100100110110;
      twice_table[1275] = 25'b1001110111000000011101000;
      twice_table[1276] = 25'b1001110110110100010011100;
      twice_table[1277] = 25'b1001110110101000001010100;
      twice_table[1278] = 25'b1001110110011100000010000;
      twice_table[1279] = 25'b1001110110001111111010000;
      twice_table[1280] = 25'b1001110110000011110010100;
      twice_table[1281] = 25'b1001110101110111101011010;
      twice_table[1282] = 25'b1001110101101011100100110;
      twice_table[1283] = 25'b1001110101011111011110100;
      twice_table[1284] = 25'b1001110101010011011000110;
      twice_table[1285] = 25'b1001110101000111010011100;
      twice_table[1286] = 25'b1001110100111011001110110;
      twice_table[1287] = 25'b1001110100101111001010100;
      twice_table[1288] = 25'b1001110100100011000110100;
      twice_table[1289] = 25'b1001110100010111000011010;
      twice_table[1290] = 25'b1001110100001011000000010;
      twice_table[1291] = 25'b1001110011111110111101110;
      twice_table[1292] = 25'b1001110011110010111011110;
      twice_table[1293] = 25'b1001110011100110111010010;
      twice_table[1294] = 25'b1001110011011010111001000;
      twice_table[1295] = 25'b1001110011001110111000100;
      twice_table[1296] = 25'b1001110011000010111000010;
      twice_table[1297] = 25'b1001110010110110111000100;
      twice_table[1298] = 25'b1001110010101010111001010;
      twice_table[1299] = 25'b1001110010011110111010100;
      twice_table[1300] = 25'b1001110010010010111100010;
      twice_table[1301] = 25'b1001110010000110111110010;
      twice_table[1302] = 25'b1001110001111011000001000;
      twice_table[1303] = 25'b1001110001101111000100000;
      twice_table[1304] = 25'b1001110001100011000111100;
      twice_table[1305] = 25'b1001110001010111001011100;
      twice_table[1306] = 25'b1001110001001011001111110;
      twice_table[1307] = 25'b1001110000111111010100110;
      twice_table[1308] = 25'b1001110000110011011010000;
      twice_table[1309] = 25'b1001110000100111011111110;
      twice_table[1310] = 25'b1001110000011011100110000;
      twice_table[1311] = 25'b1001110000001111101100110;
      twice_table[1312] = 25'b1001110000000011110011110;
      twice_table[1313] = 25'b1001101111110111111011010;
      twice_table[1314] = 25'b1001101111101100000011100;
      twice_table[1315] = 25'b1001101111100000001011110;
      twice_table[1316] = 25'b1001101111010100010100110;
      twice_table[1317] = 25'b1001101111001000011110010;
      twice_table[1318] = 25'b1001101110111100101000000;
      twice_table[1319] = 25'b1001101110110000110010010;
      twice_table[1320] = 25'b1001101110100100111101000;
      twice_table[1321] = 25'b1001101110011001001000010;
      twice_table[1322] = 25'b1001101110001101010100000;
      twice_table[1323] = 25'b1001101110000001100000000;
      twice_table[1324] = 25'b1001101101110101101100100;
      twice_table[1325] = 25'b1001101101101001111001100;
      twice_table[1326] = 25'b1001101101011110000111000;
      twice_table[1327] = 25'b1001101101010010010100110;
      twice_table[1328] = 25'b1001101101000110100011000;
      twice_table[1329] = 25'b1001101100111010110010000;
      twice_table[1330] = 25'b1001101100101111000001000;
      twice_table[1331] = 25'b1001101100100011010000110;
      twice_table[1332] = 25'b1001101100010111100001000;
      twice_table[1333] = 25'b1001101100001011110001100;
      twice_table[1334] = 25'b1001101100000000000010100;
      twice_table[1335] = 25'b1001101011110100010011110;
      twice_table[1336] = 25'b1001101011101000100101110;
      twice_table[1337] = 25'b1001101011011100111000000;
      twice_table[1338] = 25'b1001101011010001001010110;
      twice_table[1339] = 25'b1001101011000101011110000;
      twice_table[1340] = 25'b1001101010111001110001110;
      twice_table[1341] = 25'b1001101010101110000101110;
      twice_table[1342] = 25'b1001101010100010011010010;
      twice_table[1343] = 25'b1001101010010110101111010;
      twice_table[1344] = 25'b1001101010001011000100110;
      twice_table[1345] = 25'b1001101001111111011010100;
      twice_table[1346] = 25'b1001101001110011110001000;
      twice_table[1347] = 25'b1001101001101000000111100;
      twice_table[1348] = 25'b1001101001011100011110110;
      twice_table[1349] = 25'b1001101001010000110110100;
      twice_table[1350] = 25'b1001101001000101001110100;
      twice_table[1351] = 25'b1001101000111001100111000;
      twice_table[1352] = 25'b1001101000101101111111110;
      twice_table[1353] = 25'b1001101000100010011001010;
      twice_table[1354] = 25'b1001101000010110110011000;
      twice_table[1355] = 25'b1001101000001011001101010;
      twice_table[1356] = 25'b1001100111111111101000000;
      twice_table[1357] = 25'b1001100111110100000011000;
      twice_table[1358] = 25'b1001100111101000011110100;
      twice_table[1359] = 25'b1001100111011100111010100;
      twice_table[1360] = 25'b1001100111010001010111000;
      twice_table[1361] = 25'b1001100111000101110011110;
      twice_table[1362] = 25'b1001100110111010010001000;
      twice_table[1363] = 25'b1001100110101110101110110;
      twice_table[1364] = 25'b1001100110100011001101000;
      twice_table[1365] = 25'b1001100110010111101011100;
      twice_table[1366] = 25'b1001100110001100001010100;
      twice_table[1367] = 25'b1001100110000000101010000;
      twice_table[1368] = 25'b1001100101110101001001110;
      twice_table[1369] = 25'b1001100101101001101010010;
      twice_table[1370] = 25'b1001100101011110001011000;
      twice_table[1371] = 25'b1001100101010010101100000;
      twice_table[1372] = 25'b1001100101000111001101110;
      twice_table[1373] = 25'b1001100100111011101111110;
      twice_table[1374] = 25'b1001100100110000010010000;
      twice_table[1375] = 25'b1001100100100100110101000;
      twice_table[1376] = 25'b1001100100011001011000010;
      twice_table[1377] = 25'b1001100100001101111100000;
      twice_table[1378] = 25'b1001100100000010100000010;
      twice_table[1379] = 25'b1001100011110111000100110;
      twice_table[1380] = 25'b1001100011101011101001110;
      twice_table[1381] = 25'b1001100011100000001111010;
      twice_table[1382] = 25'b1001100011010100110101000;
      twice_table[1383] = 25'b1001100011001001011011100;
      twice_table[1384] = 25'b1001100010111110000010000;
      twice_table[1385] = 25'b1001100010110010101001010;
      twice_table[1386] = 25'b1001100010100111010000110;
      twice_table[1387] = 25'b1001100010011011111000110;
      twice_table[1388] = 25'b1001100010010000100001010;
      twice_table[1389] = 25'b1001100010000101001010000;
      twice_table[1390] = 25'b1001100001111001110011010;
      twice_table[1391] = 25'b1001100001101110011101000;
      twice_table[1392] = 25'b1001100001100011000111000;
      twice_table[1393] = 25'b1001100001010111110001110;
      twice_table[1394] = 25'b1001100001001100011100100;
      twice_table[1395] = 25'b1001100001000001001000000;
      twice_table[1396] = 25'b1001100000110101110011110;
      twice_table[1397] = 25'b1001100000101010100000000;
      twice_table[1398] = 25'b1001100000011111001100100;
      twice_table[1399] = 25'b1001100000010011111001110;
      twice_table[1400] = 25'b1001100000001000100111000;
      twice_table[1401] = 25'b1001011111111101010101000;
      twice_table[1402] = 25'b1001011111110010000011010;
      twice_table[1403] = 25'b1001011111100110110010000;
      twice_table[1404] = 25'b1001011111011011100001010;
      twice_table[1405] = 25'b1001011111010000010000110;
      twice_table[1406] = 25'b1001011111000101000000110;
      twice_table[1407] = 25'b1001011110111001110001010;
      twice_table[1408] = 25'b1001011110101110100010000;
      twice_table[1409] = 25'b1001011110100011010011010;
      twice_table[1410] = 25'b1001011110011000000100110;
      twice_table[1411] = 25'b1001011110001100110110110;
      twice_table[1412] = 25'b1001011110000001101001010;
      twice_table[1413] = 25'b1001011101110110011100010;
      twice_table[1414] = 25'b1001011101101011001111100;
      twice_table[1415] = 25'b1001011101100000000011010;
      twice_table[1416] = 25'b1001011101010100110111100;
      twice_table[1417] = 25'b1001011101001001101100000;
      twice_table[1418] = 25'b1001011100111110100001000;
      twice_table[1419] = 25'b1001011100110011010110010;
      twice_table[1420] = 25'b1001011100101000001100000;
      twice_table[1421] = 25'b1001011100011101000010010;
      twice_table[1422] = 25'b1001011100010001111000110;
      twice_table[1423] = 25'b1001011100000110101111110;
      twice_table[1424] = 25'b1001011011111011100111010;
      twice_table[1425] = 25'b1001011011110000011111000;
      twice_table[1426] = 25'b1001011011100101010111010;
      twice_table[1427] = 25'b1001011011011010010000000;
      twice_table[1428] = 25'b1001011011001111001001000;
      twice_table[1429] = 25'b1001011011000100000010100;
      twice_table[1430] = 25'b1001011010111000111100100;
      twice_table[1431] = 25'b1001011010101101110110110;
      twice_table[1432] = 25'b1001011010100010110001100;
      twice_table[1433] = 25'b1001011010010111101100100;
      twice_table[1434] = 25'b1001011010001100101000000;
      twice_table[1435] = 25'b1001011010000001100100000;
      twice_table[1436] = 25'b1001011001110110100000010;
      twice_table[1437] = 25'b1001011001101011011101000;
      twice_table[1438] = 25'b1001011001100000011010010;
      twice_table[1439] = 25'b1001011001010101010111110;
      twice_table[1440] = 25'b1001011001001010010101110;
      twice_table[1441] = 25'b1001011000111111010100000;
      twice_table[1442] = 25'b1001011000110100010010110;
      twice_table[1443] = 25'b1001011000101001010010000;
      twice_table[1444] = 25'b1001011000011110010001100;
      twice_table[1445] = 25'b1001011000010011010001100;
      twice_table[1446] = 25'b1001011000001000010001110;
      twice_table[1447] = 25'b1001010111111101010010100;
      twice_table[1448] = 25'b1001010111110010010011110;
      twice_table[1449] = 25'b1001010111100111010101010;
      twice_table[1450] = 25'b1001010111011100010111010;
      twice_table[1451] = 25'b1001010111010001011001110;
      twice_table[1452] = 25'b1001010111000110011100100;
      twice_table[1453] = 25'b1001010110111011011111110;
      twice_table[1454] = 25'b1001010110110000100011010;
      twice_table[1455] = 25'b1001010110100101100111010;
      twice_table[1456] = 25'b1001010110011010101011100;
      twice_table[1457] = 25'b1001010110001111110000010;
      twice_table[1458] = 25'b1001010110000100110101100;
      twice_table[1459] = 25'b1001010101111001111011010;
      twice_table[1460] = 25'b1001010101101111000001000;
      twice_table[1461] = 25'b1001010101100100000111100;
      twice_table[1462] = 25'b1001010101011001001110010;
      twice_table[1463] = 25'b1001010101001110010101100;
      twice_table[1464] = 25'b1001010101000011011101000;
      twice_table[1465] = 25'b1001010100111000100101000;
      twice_table[1466] = 25'b1001010100101101101101010;
      twice_table[1467] = 25'b1001010100100010110110000;
      twice_table[1468] = 25'b1001010100010111111111010;
      twice_table[1469] = 25'b1001010100001101001000110;
      twice_table[1470] = 25'b1001010100000010010010110;
      twice_table[1471] = 25'b1001010011110111011101000;
      twice_table[1472] = 25'b1001010011101100100111110;
      twice_table[1473] = 25'b1001010011100001110010110;
      twice_table[1474] = 25'b1001010011010110111110010;
      twice_table[1475] = 25'b1001010011001100001010010;
      twice_table[1476] = 25'b1001010011000001010110100;
      twice_table[1477] = 25'b1001010010110110100011010;
      twice_table[1478] = 25'b1001010010101011110000010;
      twice_table[1479] = 25'b1001010010100000111101110;
      twice_table[1480] = 25'b1001010010010110001011110;
      twice_table[1481] = 25'b1001010010001011011010000;
      twice_table[1482] = 25'b1001010010000000101000100;
      twice_table[1483] = 25'b1001010001110101110111110;
      twice_table[1484] = 25'b1001010001101011000111000;
      twice_table[1485] = 25'b1001010001100000010111000;
      twice_table[1486] = 25'b1001010001010101100111000;
      twice_table[1487] = 25'b1001010001001010110111110;
      twice_table[1488] = 25'b1001010001000000001000110;
      twice_table[1489] = 25'b1001010000110101011010000;
      twice_table[1490] = 25'b1001010000101010101011110;
      twice_table[1491] = 25'b1001010000011111111110000;
      twice_table[1492] = 25'b1001010000010101010000100;
      twice_table[1493] = 25'b1001010000001010100011100;
      twice_table[1494] = 25'b1001001111111111110110110;
      twice_table[1495] = 25'b1001001111110101001010100;
      twice_table[1496] = 25'b1001001111101010011110100;
      twice_table[1497] = 25'b1001001111011111110011000;
      twice_table[1498] = 25'b1001001111010101000111110;
      twice_table[1499] = 25'b1001001111001010011101000;
      twice_table[1500] = 25'b1001001110111111110010110;
      twice_table[1501] = 25'b1001001110110101001000110;
      twice_table[1502] = 25'b1001001110101010011111010;
      twice_table[1503] = 25'b1001001110011111110110000;
      twice_table[1504] = 25'b1001001110010101001101000;
      twice_table[1505] = 25'b1001001110001010100100100;
      twice_table[1506] = 25'b1001001101111111111100100;
      twice_table[1507] = 25'b1001001101110101010100110;
      twice_table[1508] = 25'b1001001101101010101101100;
      twice_table[1509] = 25'b1001001101100000000110100;
      twice_table[1510] = 25'b1001001101010101100000000;
      twice_table[1511] = 25'b1001001101001010111010000;
      twice_table[1512] = 25'b1001001101000000010100010;
      twice_table[1513] = 25'b1001001100110101101110110;
      twice_table[1514] = 25'b1001001100101011001001110;
      twice_table[1515] = 25'b1001001100100000100101000;
      twice_table[1516] = 25'b1001001100010110000000110;
      twice_table[1517] = 25'b1001001100001011011101000;
      twice_table[1518] = 25'b1001001100000000111001100;
      twice_table[1519] = 25'b1001001011110110010110010;
      twice_table[1520] = 25'b1001001011101011110011100;
      twice_table[1521] = 25'b1001001011100001010001010;
      twice_table[1522] = 25'b1001001011010110101111010;
      twice_table[1523] = 25'b1001001011001100001101100;
      twice_table[1524] = 25'b1001001011000001101100010;
      twice_table[1525] = 25'b1001001010110111001011100;
      twice_table[1526] = 25'b1001001010101100101011000;
      twice_table[1527] = 25'b1001001010100010001011000;
      twice_table[1528] = 25'b1001001010010111101011010;
      twice_table[1529] = 25'b1001001010001101001011110;
      twice_table[1530] = 25'b1001001010000010101100110;
      twice_table[1531] = 25'b1001001001111000001110010;
      twice_table[1532] = 25'b1001001001101101110000000;
      twice_table[1533] = 25'b1001001001100011010010010;
      twice_table[1534] = 25'b1001001001011000110100110;
      twice_table[1535] = 25'b1001001001001110010111100;
      twice_table[1536] = 25'b1001001001000011111010110;
      twice_table[1537] = 25'b1001001000111001011110100;
      twice_table[1538] = 25'b1001001000101111000010100;
      twice_table[1539] = 25'b1001001000100100100110110;
      twice_table[1540] = 25'b1001001000011010001011100;
      twice_table[1541] = 25'b1001001000001111110000110;
      twice_table[1542] = 25'b1001001000000101010110010;
      twice_table[1543] = 25'b1001000111111010111100000;
      twice_table[1544] = 25'b1001000111110000100010010;
      twice_table[1545] = 25'b1001000111100110001001000;
      twice_table[1546] = 25'b1001000111011011110000000;
      twice_table[1547] = 25'b1001000111010001010111010;
      twice_table[1548] = 25'b1001000111000110111111000;
      twice_table[1549] = 25'b1001000110111100100111000;
      twice_table[1550] = 25'b1001000110110010001111100;
      twice_table[1551] = 25'b1001000110100111111000100;
      twice_table[1552] = 25'b1001000110011101100001100;
      twice_table[1553] = 25'b1001000110010011001011010;
      twice_table[1554] = 25'b1001000110001000110101000;
      twice_table[1555] = 25'b1001000101111110011111100;
      twice_table[1556] = 25'b1001000101110100001010000;
      twice_table[1557] = 25'b1001000101101001110101000;
      twice_table[1558] = 25'b1001000101011111100000100;
      twice_table[1559] = 25'b1001000101010101001100010;
      twice_table[1560] = 25'b1001000101001010111000100;
      twice_table[1561] = 25'b1001000101000000100101000;
      twice_table[1562] = 25'b1001000100110110010001110;
      twice_table[1563] = 25'b1001000100101011111111000;
      twice_table[1564] = 25'b1001000100100001101100100;
      twice_table[1565] = 25'b1001000100010111011010100;
      twice_table[1566] = 25'b1001000100001101001000110;
      twice_table[1567] = 25'b1001000100000010110111100;
      twice_table[1568] = 25'b1001000011111000100110100;
      twice_table[1569] = 25'b1001000011101110010110000;
      twice_table[1570] = 25'b1001000011100100000101110;
      twice_table[1571] = 25'b1001000011011001110110000;
      twice_table[1572] = 25'b1001000011001111100110100;
      twice_table[1573] = 25'b1001000011000101010111010;
      twice_table[1574] = 25'b1001000010111011001000100;
      twice_table[1575] = 25'b1001000010110000111010000;
      twice_table[1576] = 25'b1001000010100110101100000;
      twice_table[1577] = 25'b1001000010011100011110010;
      twice_table[1578] = 25'b1001000010010010010001000;
      twice_table[1579] = 25'b1001000010001000000100000;
      twice_table[1580] = 25'b1001000001111101110111100;
      twice_table[1581] = 25'b1001000001110011101011010;
      twice_table[1582] = 25'b1001000001101001011111010;
      twice_table[1583] = 25'b1001000001011111010011110;
      twice_table[1584] = 25'b1001000001010101001000100;
      twice_table[1585] = 25'b1001000001001010111101110;
      twice_table[1586] = 25'b1001000001000000110011010;
      twice_table[1587] = 25'b1001000000110110101001010;
      twice_table[1588] = 25'b1001000000101100011111100;
      twice_table[1589] = 25'b1001000000100010010110000;
      twice_table[1590] = 25'b1001000000011000001101000;
      twice_table[1591] = 25'b1001000000001110000100010;
      twice_table[1592] = 25'b1001000000000011111100000;
      twice_table[1593] = 25'b1000111111111001110100000;
      twice_table[1594] = 25'b1000111111101111101100100;
      twice_table[1595] = 25'b1000111111100101100101010;
      twice_table[1596] = 25'b1000111111011011011110010;
      twice_table[1597] = 25'b1000111111010001010111110;
      twice_table[1598] = 25'b1000111111000111010001100;
      twice_table[1599] = 25'b1000111110111101001011110;
      twice_table[1600] = 25'b1000111110110011000110010;
      twice_table[1601] = 25'b1000111110101001000001010;
      twice_table[1602] = 25'b1000111110011110111100100;
      twice_table[1603] = 25'b1000111110010100111000000;
      twice_table[1604] = 25'b1000111110001010110100000;
      twice_table[1605] = 25'b1000111110000000110000010;
      twice_table[1606] = 25'b1000111101110110101100110;
      twice_table[1607] = 25'b1000111101101100101001110;
      twice_table[1608] = 25'b1000111101100010100111010;
      twice_table[1609] = 25'b1000111101011000100101000;
      twice_table[1610] = 25'b1000111101001110100011000;
      twice_table[1611] = 25'b1000111101000100100001010;
      twice_table[1612] = 25'b1000111100111010100000000;
      twice_table[1613] = 25'b1000111100110000011111010;
      twice_table[1614] = 25'b1000111100100110011110110;
      twice_table[1615] = 25'b1000111100011100011110100;
      twice_table[1616] = 25'b1000111100010010011110100;
      twice_table[1617] = 25'b1000111100001000011111000;
      twice_table[1618] = 25'b1000111011111110100000000;
      twice_table[1619] = 25'b1000111011110100100001000;
      twice_table[1620] = 25'b1000111011101010100010110;
      twice_table[1621] = 25'b1000111011100000100100100;
      twice_table[1622] = 25'b1000111011010110100110110;
      twice_table[1623] = 25'b1000111011001100101001100;
      twice_table[1624] = 25'b1000111011000010101100010;
      twice_table[1625] = 25'b1000111010111000101111100;
      twice_table[1626] = 25'b1000111010101110110011010;
      twice_table[1627] = 25'b1000111010100100110111010;
      twice_table[1628] = 25'b1000111010011010111011100;
      twice_table[1629] = 25'b1000111010010001000000010;
      twice_table[1630] = 25'b1000111010000111000101010;
      twice_table[1631] = 25'b1000111001111101001010100;
      twice_table[1632] = 25'b1000111001110011010000010;
      twice_table[1633] = 25'b1000111001101001010110010;
      twice_table[1634] = 25'b1000111001011111011100110;
      twice_table[1635] = 25'b1000111001010101100011100;
      twice_table[1636] = 25'b1000111001001011101010100;
      twice_table[1637] = 25'b1000111001000001110010000;
      twice_table[1638] = 25'b1000111000110111111001110;
      twice_table[1639] = 25'b1000111000101110000001110;
      twice_table[1640] = 25'b1000111000100100001010010;
      twice_table[1641] = 25'b1000111000011010010011000;
      twice_table[1642] = 25'b1000111000010000011100010;
      twice_table[1643] = 25'b1000111000000110100101110;
      twice_table[1644] = 25'b1000110111111100101111100;
      twice_table[1645] = 25'b1000110111110010111001100;
      twice_table[1646] = 25'b1000110111101001000100000;
      twice_table[1647] = 25'b1000110111011111001111000;
      twice_table[1648] = 25'b1000110111010101011010010;
      twice_table[1649] = 25'b1000110111001011100101110;
      twice_table[1650] = 25'b1000110111000001110001100;
      twice_table[1651] = 25'b1000110110110111111101110;
      twice_table[1652] = 25'b1000110110101110001010010;
      twice_table[1653] = 25'b1000110110100100010111010;
      twice_table[1654] = 25'b1000110110011010100100010;
      twice_table[1655] = 25'b1000110110010000110010000;
      twice_table[1656] = 25'b1000110110000110111111110;
      twice_table[1657] = 25'b1000110101111101001110000;
      twice_table[1658] = 25'b1000110101110011011100100;
      twice_table[1659] = 25'b1000110101101001101011100;
      twice_table[1660] = 25'b1000110101011111111010110;
      twice_table[1661] = 25'b1000110101010110001010010;
      twice_table[1662] = 25'b1000110101001100011010010;
      twice_table[1663] = 25'b1000110101000010101010100;
      twice_table[1664] = 25'b1000110100111000111011000;
      twice_table[1665] = 25'b1000110100101111001100000;
      twice_table[1666] = 25'b1000110100100101011101010;
      twice_table[1667] = 25'b1000110100011011101111000;
      twice_table[1668] = 25'b1000110100010010000000110;
      twice_table[1669] = 25'b1000110100001000010011000;
      twice_table[1670] = 25'b1000110011111110100101110;
      twice_table[1671] = 25'b1000110011110100111000100;
      twice_table[1672] = 25'b1000110011101011001100000;
      twice_table[1673] = 25'b1000110011100001011111100;
      twice_table[1674] = 25'b1000110011010111110011100;
      twice_table[1675] = 25'b1000110011001110000111110;
      twice_table[1676] = 25'b1000110011000100011100010;
      twice_table[1677] = 25'b1000110010111010110001010;
      twice_table[1678] = 25'b1000110010110001000110100;
      twice_table[1679] = 25'b1000110010100111011100000;
      twice_table[1680] = 25'b1000110010011101110010000;
      twice_table[1681] = 25'b1000110010010100001000010;
      twice_table[1682] = 25'b1000110010001010011110110;
      twice_table[1683] = 25'b1000110010000000110101110;
      twice_table[1684] = 25'b1000110001110111001101000;
      twice_table[1685] = 25'b1000110001101101100100100;
      twice_table[1686] = 25'b1000110001100011111100100;
      twice_table[1687] = 25'b1000110001011010010100110;
      twice_table[1688] = 25'b1000110001010000101101010;
      twice_table[1689] = 25'b1000110001000111000110010;
      twice_table[1690] = 25'b1000110000111101011111100;
      twice_table[1691] = 25'b1000110000110011111001000;
      twice_table[1692] = 25'b1000110000101010010011000;
      twice_table[1693] = 25'b1000110000100000101101010;
      twice_table[1694] = 25'b1000110000010111000111110;
      twice_table[1695] = 25'b1000110000001101100010100;
      twice_table[1696] = 25'b1000110000000011111101110;
      twice_table[1697] = 25'b1000101111111010011001010;
      twice_table[1698] = 25'b1000101111110000110101010;
      twice_table[1699] = 25'b1000101111100111010001010;
      twice_table[1700] = 25'b1000101111011101101101110;
      twice_table[1701] = 25'b1000101111010100001010110;
      twice_table[1702] = 25'b1000101111001010100111110;
      twice_table[1703] = 25'b1000101111000001000101010;
      twice_table[1704] = 25'b1000101110110111100011010;
      twice_table[1705] = 25'b1000101110101110000001010;
      twice_table[1706] = 25'b1000101110100100011111110;
      twice_table[1707] = 25'b1000101110011010111110100;
      twice_table[1708] = 25'b1000101110010001011101110;
      twice_table[1709] = 25'b1000101110000111111101000;
      twice_table[1710] = 25'b1000101101111110011100110;
      twice_table[1711] = 25'b1000101101110100111101000;
      twice_table[1712] = 25'b1000101101101011011101010;
      twice_table[1713] = 25'b1000101101100001111110000;
      twice_table[1714] = 25'b1000101101011000011111000;
      twice_table[1715] = 25'b1000101101001111000000100;
      twice_table[1716] = 25'b1000101101000101100010010;
      twice_table[1717] = 25'b1000101100111100000100010;
      twice_table[1718] = 25'b1000101100110010100110100;
      twice_table[1719] = 25'b1000101100101001001001010;
      twice_table[1720] = 25'b1000101100011111101100010;
      twice_table[1721] = 25'b1000101100010110001111100;
      twice_table[1722] = 25'b1000101100001100110011000;
      twice_table[1723] = 25'b1000101100000011010111000;
      twice_table[1724] = 25'b1000101011111001111011010;
      twice_table[1725] = 25'b1000101011110000100000000;
      twice_table[1726] = 25'b1000101011100111000100110;
      twice_table[1727] = 25'b1000101011011101101010000;
      twice_table[1728] = 25'b1000101011010100001111100;
      twice_table[1729] = 25'b1000101011001010110101100;
      twice_table[1730] = 25'b1000101011000001011011100;
      twice_table[1731] = 25'b1000101010111000000010000;
      twice_table[1732] = 25'b1000101010101110101001000;
      twice_table[1733] = 25'b1000101010100101010000000;
      twice_table[1734] = 25'b1000101010011011110111100;
      twice_table[1735] = 25'b1000101010010010011111010;
      twice_table[1736] = 25'b1000101010001001000111010;
      twice_table[1737] = 25'b1000101001111111101111110;
      twice_table[1738] = 25'b1000101001110110011000100;
      twice_table[1739] = 25'b1000101001101101000001100;
      twice_table[1740] = 25'b1000101001100011101011000;
      twice_table[1741] = 25'b1000101001011010010100100;
      twice_table[1742] = 25'b1000101001010000111110100;
      twice_table[1743] = 25'b1000101001000111101000110;
      twice_table[1744] = 25'b1000101000111110010011100;
      twice_table[1745] = 25'b1000101000110100111110100;
      twice_table[1746] = 25'b1000101000101011101001110;
      twice_table[1747] = 25'b1000101000100010010101010;
      twice_table[1748] = 25'b1000101000011001000001000;
      twice_table[1749] = 25'b1000101000001111101101010;
      twice_table[1750] = 25'b1000101000000110011001110;
      twice_table[1751] = 25'b1000100111111101000110100;
      twice_table[1752] = 25'b1000100111110011110011110;
      twice_table[1753] = 25'b1000100111101010100001010;
      twice_table[1754] = 25'b1000100111100001001111000;
      twice_table[1755] = 25'b1000100111010111111101000;
      twice_table[1756] = 25'b1000100111001110101011010;
      twice_table[1757] = 25'b1000100111000101011010000;
      twice_table[1758] = 25'b1000100110111100001001000;
      twice_table[1759] = 25'b1000100110110010111000010;
      twice_table[1760] = 25'b1000100110101001101000000;
      twice_table[1761] = 25'b1000100110100000011000000;
      twice_table[1762] = 25'b1000100110010111001000010;
      twice_table[1763] = 25'b1000100110001101111000110;
      twice_table[1764] = 25'b1000100110000100101001100;
      twice_table[1765] = 25'b1000100101111011011010110;
      twice_table[1766] = 25'b1000100101110010001100010;
      twice_table[1767] = 25'b1000100101101000111110000;
      twice_table[1768] = 25'b1000100101011111110000010;
      twice_table[1769] = 25'b1000100101010110100010100;
      twice_table[1770] = 25'b1000100101001101010101010;
      twice_table[1771] = 25'b1000100101000100001000010;
      twice_table[1772] = 25'b1000100100111010111011110;
      twice_table[1773] = 25'b1000100100110001101111010;
      twice_table[1774] = 25'b1000100100101000100011010;
      twice_table[1775] = 25'b1000100100011111010111100;
      twice_table[1776] = 25'b1000100100010110001100010;
      twice_table[1777] = 25'b1000100100001101000001000;
      twice_table[1778] = 25'b1000100100000011110110010;
      twice_table[1779] = 25'b1000100011111010101011110;
      twice_table[1780] = 25'b1000100011110001100001100;
      twice_table[1781] = 25'b1000100011101000010111100;
      twice_table[1782] = 25'b1000100011011111001110000;
      twice_table[1783] = 25'b1000100011010110000100110;
      twice_table[1784] = 25'b1000100011001100111011110;
      twice_table[1785] = 25'b1000100011000011110011000;
      twice_table[1786] = 25'b1000100010111010101010110;
      twice_table[1787] = 25'b1000100010110001100010110;
      twice_table[1788] = 25'b1000100010101000011011000;
      twice_table[1789] = 25'b1000100010011111010011100;
      twice_table[1790] = 25'b1000100010010110001100010;
      twice_table[1791] = 25'b1000100010001101000101100;
      twice_table[1792] = 25'b1000100010000011111111000;
      twice_table[1793] = 25'b1000100001111010111000110;
      twice_table[1794] = 25'b1000100001110001110010110;
      twice_table[1795] = 25'b1000100001101000101101000;
      twice_table[1796] = 25'b1000100001011111100111110;
      twice_table[1797] = 25'b1000100001010110100010110;
      twice_table[1798] = 25'b1000100001001101011110000;
      twice_table[1799] = 25'b1000100001000100011001100;
      twice_table[1800] = 25'b1000100000111011010101100;
      twice_table[1801] = 25'b1000100000110010010001110;
      twice_table[1802] = 25'b1000100000101001001110000;
      twice_table[1803] = 25'b1000100000100000001011000;
      twice_table[1804] = 25'b1000100000010111001000000;
      twice_table[1805] = 25'b1000100000001110000101010;
      twice_table[1806] = 25'b1000100000000101000011000;
      twice_table[1807] = 25'b1000011111111100000001000;
      twice_table[1808] = 25'b1000011111110010111111010;
      twice_table[1809] = 25'b1000011111101001111110000;
      twice_table[1810] = 25'b1000011111100000111100110;
      twice_table[1811] = 25'b1000011111010111111100000;
      twice_table[1812] = 25'b1000011111001110111011100;
      twice_table[1813] = 25'b1000011111000101111011010;
      twice_table[1814] = 25'b1000011110111100111011010;
      twice_table[1815] = 25'b1000011110110011111011110;
      twice_table[1816] = 25'b1000011110101010111100010;
      twice_table[1817] = 25'b1000011110100001111101010;
      twice_table[1818] = 25'b1000011110011000111110100;
      twice_table[1819] = 25'b1000011110010000000000010;
      twice_table[1820] = 25'b1000011110000111000010000;
      twice_table[1821] = 25'b1000011101111110000100010;
      twice_table[1822] = 25'b1000011101110101000110100;
      twice_table[1823] = 25'b1000011101101100001001010;
      twice_table[1824] = 25'b1000011101100011001100100;
      twice_table[1825] = 25'b1000011101011010001111110;
      twice_table[1826] = 25'b1000011101010001010011100;
      twice_table[1827] = 25'b1000011101001000010111010;
      twice_table[1828] = 25'b1000011100111111011011100;
      twice_table[1829] = 25'b1000011100110110100000000;
      twice_table[1830] = 25'b1000011100101101100101000;
      twice_table[1831] = 25'b1000011100100100101010000;
      twice_table[1832] = 25'b1000011100011011101111100;
      twice_table[1833] = 25'b1000011100010010110101000;
      twice_table[1834] = 25'b1000011100001001111011000;
      twice_table[1835] = 25'b1000011100000001000001100;
      twice_table[1836] = 25'b1000011011111000001000000;
      twice_table[1837] = 25'b1000011011101111001110110;
      twice_table[1838] = 25'b1000011011100110010110000;
      twice_table[1839] = 25'b1000011011011101011101100;
      twice_table[1840] = 25'b1000011011010100100101010;
      twice_table[1841] = 25'b1000011011001011101101010;
      twice_table[1842] = 25'b1000011011000010110101100;
      twice_table[1843] = 25'b1000011010111001111110010;
      twice_table[1844] = 25'b1000011010110001000111010;
      twice_table[1845] = 25'b1000011010101000010000010;
      twice_table[1846] = 25'b1000011010011111011001110;
      twice_table[1847] = 25'b1000011010010110100011110;
      twice_table[1848] = 25'b1000011010001101101101110;
      twice_table[1849] = 25'b1000011010000100111000010;
      twice_table[1850] = 25'b1000011001111100000010110;
      twice_table[1851] = 25'b1000011001110011001101110;
      twice_table[1852] = 25'b1000011001101010011001000;
      twice_table[1853] = 25'b1000011001100001100100100;
      twice_table[1854] = 25'b1000011001011000110000010;
      twice_table[1855] = 25'b1000011001001111111100100;
      twice_table[1856] = 25'b1000011001000111001000110;
      twice_table[1857] = 25'b1000011000111110010101100;
      twice_table[1858] = 25'b1000011000110101100010100;
      twice_table[1859] = 25'b1000011000101100101111110;
      twice_table[1860] = 25'b1000011000100011111101010;
      twice_table[1861] = 25'b1000011000011011001011010;
      twice_table[1862] = 25'b1000011000010010011001010;
      twice_table[1863] = 25'b1000011000001001100111110;
      twice_table[1864] = 25'b1000011000000000110110100;
      twice_table[1865] = 25'b1000010111111000000101100;
      twice_table[1866] = 25'b1000010111101111010100110;
      twice_table[1867] = 25'b1000010111100110100100010;
      twice_table[1868] = 25'b1000010111011101110100000;
      twice_table[1869] = 25'b1000010111010101000100010;
      twice_table[1870] = 25'b1000010111001100010100110;
      twice_table[1871] = 25'b1000010111000011100101100;
      twice_table[1872] = 25'b1000010110111010110110100;
      twice_table[1873] = 25'b1000010110110010000111110;
      twice_table[1874] = 25'b1000010110101001011001010;
      twice_table[1875] = 25'b1000010110100000101011000;
      twice_table[1876] = 25'b1000010110010111111101010;
      twice_table[1877] = 25'b1000010110001111001111100;
      twice_table[1878] = 25'b1000010110000110100010010;
      twice_table[1879] = 25'b1000010101111101110101010;
      twice_table[1880] = 25'b1000010101110101001000100;
      twice_table[1881] = 25'b1000010101101100011100000;
      twice_table[1882] = 25'b1000010101100011110000000;
      twice_table[1883] = 25'b1000010101011011000100000;
      twice_table[1884] = 25'b1000010101010010011000100;
      twice_table[1885] = 25'b1000010101001001101101010;
      twice_table[1886] = 25'b1000010101000001000010000;
      twice_table[1887] = 25'b1000010100111000010111010;
      twice_table[1888] = 25'b1000010100101111101101000;
      twice_table[1889] = 25'b1000010100100111000010110;
      twice_table[1890] = 25'b1000010100011110011000110;
      twice_table[1891] = 25'b1000010100010101101111010;
      twice_table[1892] = 25'b1000010100001101000101110;
      twice_table[1893] = 25'b1000010100000100011100110;
      twice_table[1894] = 25'b1000010011111011110100000;
      twice_table[1895] = 25'b1000010011110011001011100;
      twice_table[1896] = 25'b1000010011101010100011010;
      twice_table[1897] = 25'b1000010011100001111011010;
      twice_table[1898] = 25'b1000010011011001010011100;
      twice_table[1899] = 25'b1000010011010000101100010;
      twice_table[1900] = 25'b1000010011001000000101000;
      twice_table[1901] = 25'b1000010010111111011110010;
      twice_table[1902] = 25'b1000010010110110110111110;
      twice_table[1903] = 25'b1000010010101110010001100;
      twice_table[1904] = 25'b1000010010100101101011100;
      twice_table[1905] = 25'b1000010010011101000101110;
      twice_table[1906] = 25'b1000010010010100100000010;
      twice_table[1907] = 25'b1000010010001011111011010;
      twice_table[1908] = 25'b1000010010000011010110010;
      twice_table[1909] = 25'b1000010001111010110001110;
      twice_table[1910] = 25'b1000010001110010001101010;
      twice_table[1911] = 25'b1000010001101001101001010;
      twice_table[1912] = 25'b1000010001100001000101100;
      twice_table[1913] = 25'b1000010001011000100010000;
      twice_table[1914] = 25'b1000010001001111111110110;
      twice_table[1915] = 25'b1000010001000111011100000;
      twice_table[1916] = 25'b1000010000111110111001010;
      twice_table[1917] = 25'b1000010000110110010110110;
      twice_table[1918] = 25'b1000010000101101110100110;
      twice_table[1919] = 25'b1000010000100101010011000;
      twice_table[1920] = 25'b1000010000011100110001010;
      twice_table[1921] = 25'b1000010000010100010000000;
      twice_table[1922] = 25'b1000010000001011101111000;
      twice_table[1923] = 25'b1000010000000011001110010;
      twice_table[1924] = 25'b1000001111111010101101110;
      twice_table[1925] = 25'b1000001111110010001101100;
      twice_table[1926] = 25'b1000001111101001101101110;
      twice_table[1927] = 25'b1000001111100001001110000;
      twice_table[1928] = 25'b1000001111011000101110110;
      twice_table[1929] = 25'b1000001111010000001111100;
      twice_table[1930] = 25'b1000001111000111110000110;
      twice_table[1931] = 25'b1000001110111111010010010;
      twice_table[1932] = 25'b1000001110110110110100000;
      twice_table[1933] = 25'b1000001110101110010110000;
      twice_table[1934] = 25'b1000001110100101111000010;
      twice_table[1935] = 25'b1000001110011101011010110;
      twice_table[1936] = 25'b1000001110010100111101100;
      twice_table[1937] = 25'b1000001110001100100000100;
      twice_table[1938] = 25'b1000001110000100000100000;
      twice_table[1939] = 25'b1000001101111011100111100;
      twice_table[1940] = 25'b1000001101110011001011100;
      twice_table[1941] = 25'b1000001101101010101111110;
      twice_table[1942] = 25'b1000001101100010010100000;
      twice_table[1943] = 25'b1000001101011001111000110;
      twice_table[1944] = 25'b1000001101010001011101110;
      twice_table[1945] = 25'b1000001101001001000011000;
      twice_table[1946] = 25'b1000001101000000101000100;
      twice_table[1947] = 25'b1000001100111000001110010;
      twice_table[1948] = 25'b1000001100101111110100010;
      twice_table[1949] = 25'b1000001100100111011010110;
      twice_table[1950] = 25'b1000001100011111000001010;
      twice_table[1951] = 25'b1000001100010110101000000;
      twice_table[1952] = 25'b1000001100001110001111010;
      twice_table[1953] = 25'b1000001100000101110110110;
      twice_table[1954] = 25'b1000001011111101011110010;
      twice_table[1955] = 25'b1000001011110101000110010;
      twice_table[1956] = 25'b1000001011101100101110100;
      twice_table[1957] = 25'b1000001011100100010111000;
      twice_table[1958] = 25'b1000001011011011111111110;
      twice_table[1959] = 25'b1000001011010011101000110;
      twice_table[1960] = 25'b1000001011001011010010000;
      twice_table[1961] = 25'b1000001011000010111011100;
      twice_table[1962] = 25'b1000001010111010100101010;
      twice_table[1963] = 25'b1000001010110010001111010;
      twice_table[1964] = 25'b1000001010101001111001110;
      twice_table[1965] = 25'b1000001010100001100100010;
      twice_table[1966] = 25'b1000001010011001001111010;
      twice_table[1967] = 25'b1000001010010000111010010;
      twice_table[1968] = 25'b1000001010001000100101110;
      twice_table[1969] = 25'b1000001010000000010001010;
      twice_table[1970] = 25'b1000001001110111111101010;
      twice_table[1971] = 25'b1000001001101111101001100;
      twice_table[1972] = 25'b1000001001100111010110000;
      twice_table[1973] = 25'b1000001001011111000010110;
      twice_table[1974] = 25'b1000001001010110101111100;
      twice_table[1975] = 25'b1000001001001110011100110;
      twice_table[1976] = 25'b1000001001000110001010100;
      twice_table[1977] = 25'b1000001000111101111000010;
      twice_table[1978] = 25'b1000001000110101100110010;
      twice_table[1979] = 25'b1000001000101101010100100;
      twice_table[1980] = 25'b1000001000100101000011000;
      twice_table[1981] = 25'b1000001000011100110010000;
      twice_table[1982] = 25'b1000001000010100100001000;
      twice_table[1983] = 25'b1000001000001100010000010;
      twice_table[1984] = 25'b1000001000000100000000000;
      twice_table[1985] = 25'b1000000111111011101111110;
      twice_table[1986] = 25'b1000000111110011100000000;
      twice_table[1987] = 25'b1000000111101011010000100;
      twice_table[1988] = 25'b1000000111100011000001000;
      twice_table[1989] = 25'b1000000111011010110010000;
      twice_table[1990] = 25'b1000000111010010100011010;
      twice_table[1991] = 25'b1000000111001010010100100;
      twice_table[1992] = 25'b1000000111000010000110010;
      twice_table[1993] = 25'b1000000110111001111000010;
      twice_table[1994] = 25'b1000000110110001101010100;
      twice_table[1995] = 25'b1000000110101001011101000;
      twice_table[1996] = 25'b1000000110100001001111110;
      twice_table[1997] = 25'b1000000110011001000010110;
      twice_table[1998] = 25'b1000000110010000110110000;
      twice_table[1999] = 25'b1000000110001000101001100;
      twice_table[2000] = 25'b1000000110000000011101010;
      twice_table[2001] = 25'b1000000101111000010001100;
      twice_table[2002] = 25'b1000000101110000000101110;
      twice_table[2003] = 25'b1000000101100111111010010;
      twice_table[2004] = 25'b1000000101011111101111000;
      twice_table[2005] = 25'b1000000101010111100100010;
      twice_table[2006] = 25'b1000000101001111011001100;
      twice_table[2007] = 25'b1000000101000111001111000;
      twice_table[2008] = 25'b1000000100111111000101000;
      twice_table[2009] = 25'b1000000100110110111011000;
      twice_table[2010] = 25'b1000000100101110110001100;
      twice_table[2011] = 25'b1000000100100110101000000;
      twice_table[2012] = 25'b1000000100011110011111000;
      twice_table[2013] = 25'b1000000100010110010110000;
      twice_table[2014] = 25'b1000000100001110001101100;
      twice_table[2015] = 25'b1000000100000110000101000;
      twice_table[2016] = 25'b1000000011111101111101000;
      twice_table[2017] = 25'b1000000011110101110101010;
      twice_table[2018] = 25'b1000000011101101101101100;
      twice_table[2019] = 25'b1000000011100101100110010;
      twice_table[2020] = 25'b1000000011011101011111010;
      twice_table[2021] = 25'b1000000011010101011000010;
      twice_table[2022] = 25'b1000000011001101010001110;
      twice_table[2023] = 25'b1000000011000101001011100;
      twice_table[2024] = 25'b1000000010111101000101100;
      twice_table[2025] = 25'b1000000010110100111111110;
      twice_table[2026] = 25'b1000000010101100111010000;
      twice_table[2027] = 25'b1000000010100100110100110;
      twice_table[2028] = 25'b1000000010011100101111110;
      twice_table[2029] = 25'b1000000010010100101011000;
      twice_table[2030] = 25'b1000000010001100100110100;
      twice_table[2031] = 25'b1000000010000100100010010;
      twice_table[2032] = 25'b1000000001111100011110010;
      twice_table[2033] = 25'b1000000001110100011010010;
      twice_table[2034] = 25'b1000000001101100010110110;
      twice_table[2035] = 25'b1000000001100100010011100;
      twice_table[2036] = 25'b1000000001011100010000100;
      twice_table[2037] = 25'b1000000001010100001101110;
      twice_table[2038] = 25'b1000000001001100001011010;
      twice_table[2039] = 25'b1000000001000100001001000;
      twice_table[2040] = 25'b1000000000111100000111000;
      twice_table[2041] = 25'b1000000000110100000101010;
      twice_table[2042] = 25'b1000000000101100000011110;
      twice_table[2043] = 25'b1000000000100100000010100;
      twice_table[2044] = 25'b1000000000011100000001100;
      twice_table[2045] = 25'b1000000000010100000000110;
      twice_table[2046] = 25'b1000000000001100000000010;
      twice_table[2047] = 25'b1000000000000100000000000;

      square_table[0] = 25'b0111111111110000000000011;
      square_table[1] = 25'b0111111111010000000011011;
      square_table[2] = 25'b0111111110110000001001011;
      square_table[3] = 25'b0111111110010000010010011;
      square_table[4] = 25'b0111111101110000011110011;
      square_table[5] = 25'b0111111101010000101101010;
      square_table[6] = 25'b0111111100110000111111000;
      square_table[7] = 25'b0111111100010001010011111;
      square_table[8] = 25'b0111111011110001101011111;
      square_table[9] = 25'b0111111011010010000110100;
      square_table[10] = 25'b0111111010110010100100011;
      square_table[11] = 25'b0111111010010011000100111;
      square_table[12] = 25'b0111111001110011101000011;
      square_table[13] = 25'b0111111001010100001110111;
      square_table[14] = 25'b0111111000110100111000011;
      square_table[15] = 25'b0111111000010101100100111;
      square_table[16] = 25'b0111110111110110010100000;
      square_table[17] = 25'b0111110111010111000110010;
      square_table[18] = 25'b0111110110110111111011011;
      square_table[19] = 25'b0111110110011000110011010;
      square_table[20] = 25'b0111110101111001101110000;
      square_table[21] = 25'b0111110101011010101011111;
      square_table[22] = 25'b0111110100111011101100011;
      square_table[23] = 25'b0111110100011100101111111;
      square_table[24] = 25'b0111110011111101110110011;
      square_table[25] = 25'b0111110011011110111111011;
      square_table[26] = 25'b0111110011000000001011100;
      square_table[27] = 25'b0111110010100001011010011;
      square_table[28] = 25'b0111110010000010101100000;
      square_table[29] = 25'b0111110001100100000000111;
      square_table[30] = 25'b0111110001000101011000001;
      square_table[31] = 25'b0111110000100110110010100;
      square_table[32] = 25'b0111110000001000001111100;
      square_table[33] = 25'b0111101111101001101111100;
      square_table[34] = 25'b0111101111001011010010001;
      square_table[35] = 25'b0111101110101100110111101;
      square_table[36] = 25'b0111101110001110100000000;
      square_table[37] = 25'b0111101101110000001011001;
      square_table[38] = 25'b0111101101010001111001000;
      square_table[39] = 25'b0111101100110011101001101;
      square_table[40] = 25'b0111101100010101011101001;
      square_table[41] = 25'b0111101011110111010011010;
      square_table[42] = 25'b0111101011011001001100010;
      square_table[43] = 25'b0111101010111011001000001;
      square_table[44] = 25'b0111101010011101000110110;
      square_table[45] = 25'b0111101001111111000111111;
      square_table[46] = 25'b0111101001100001001011111;
      square_table[47] = 25'b0111101001000011010010101;
      square_table[48] = 25'b0111101000100101011100001;
      square_table[49] = 25'b0111101000000111101000100;
      square_table[50] = 25'b0111100111101001110111100;
      square_table[51] = 25'b0111100111001100001001001;
      square_table[52] = 25'b0111100110101110011101011;
      square_table[53] = 25'b0111100110010000110100101;
      square_table[54] = 25'b0111100101110011001110011;
      square_table[55] = 25'b0111100101010101101010111;
      square_table[56] = 25'b0111100100111000001010001;
      square_table[57] = 25'b0111100100011010101100001;
      square_table[58] = 25'b0111100011111101010000101;
      square_table[59] = 25'b0111100011011111110111111;
      square_table[60] = 25'b0111100011000010100001111;
      square_table[61] = 25'b0111100010100101001110100;
      square_table[62] = 25'b0111100010000111111101101;
      square_table[63] = 25'b0111100001101010101111101;
      square_table[64] = 25'b0111100001001101100100010;
      square_table[65] = 25'b0111100000110000011011100;
      square_table[66] = 25'b0111100000010011010101100;
      square_table[67] = 25'b0111011111110110010001111;
      square_table[68] = 25'b0111011111011001010001010;
      square_table[69] = 25'b0111011110111100010011000;
      square_table[70] = 25'b0111011110011111010111010;
      square_table[71] = 25'b0111011110000010011110011;
      square_table[72] = 25'b0111011101100101101000000;
      square_table[73] = 25'b0111011101001000110100010;
      square_table[74] = 25'b0111011100101100000011010;
      square_table[75] = 25'b0111011100001111010100100;
      square_table[76] = 25'b0111011011110010101000110;
      square_table[77] = 25'b0111011011010101111111011;
      square_table[78] = 25'b0111011010111001011000101;
      square_table[79] = 25'b0111011010011100110100011;
      square_table[80] = 25'b0111011010000000010010111;
      square_table[81] = 25'b0111011001100011110011110;
      square_table[82] = 25'b0111011001000111010111011;
      square_table[83] = 25'b0111011000101010111101011;
      square_table[84] = 25'b0111011000001110100110000;
      square_table[85] = 25'b0111010111110010010001010;
      square_table[86] = 25'b0111010111010101111111000;
      square_table[87] = 25'b0111010110111001101111011;
      square_table[88] = 25'b0111010110011101100010001;
      square_table[89] = 25'b0111010110000001010111100;
      square_table[90] = 25'b0111010101100101001111101;
      square_table[91] = 25'b0111010101001001001010000;
      square_table[92] = 25'b0111010100101101000110111;
      square_table[93] = 25'b0111010100010001000110010;
      square_table[94] = 25'b0111010011110101001000001;
      square_table[95] = 25'b0111010011011001001100111;
      square_table[96] = 25'b0111010010111101010011110;
      square_table[97] = 25'b0111010010100001011101010;
      square_table[98] = 25'b0111010010000101101001001;
      square_table[99] = 25'b0111010001101001110111100;
      square_table[100] = 25'b0111010001001110001000100;
      square_table[101] = 25'b0111010000110010011011111;
      square_table[102] = 25'b0111010000010110110001110;
      square_table[103] = 25'b0111001111111011001010010;
      square_table[104] = 25'b0111001111011111100100111;
      square_table[105] = 25'b0111001111000100000010010;
      square_table[106] = 25'b0111001110101000100001111;
      square_table[107] = 25'b0111001110001101000100001;
      square_table[108] = 25'b0111001101110001101000110;
      square_table[109] = 25'b0111001101010110001111110;
      square_table[110] = 25'b0111001100111010111001010;
      square_table[111] = 25'b0111001100011111100101000;
      square_table[112] = 25'b0111001100000100010011100;
      square_table[113] = 25'b0111001011101001000100010;
      square_table[114] = 25'b0111001011001101110111011;
      square_table[115] = 25'b0111001010110010101101000;
      square_table[116] = 25'b0111001010010111100101000;
      square_table[117] = 25'b0111001001111100011111011;
      square_table[118] = 25'b0111001001100001011100011;
      square_table[119] = 25'b0111001001000110011011100;
      square_table[120] = 25'b0111001000101011011101001;
      square_table[121] = 25'b0111001000010000100001000;
      square_table[122] = 25'b0111000111110101100111011;
      square_table[123] = 25'b0111000111011010110000001;
      square_table[124] = 25'b0111000110111111111011010;
      square_table[125] = 25'b0111000110100101001000110;
      square_table[126] = 25'b0111000110001010011000100;
      square_table[127] = 25'b0111000101101111101010110;
      square_table[128] = 25'b0111000101010100111111010;
      square_table[129] = 25'b0111000100111010010110011;
      square_table[130] = 25'b0111000100011111101111100;
      square_table[131] = 25'b0111000100000101001011010;
      square_table[132] = 25'b0111000011101010101001010;
      square_table[133] = 25'b0111000011010000001001011;
      square_table[134] = 25'b0111000010110101101100001;
      square_table[135] = 25'b0111000010011011010001001;
      square_table[136] = 25'b0111000010000000111000010;
      square_table[137] = 25'b0111000001100110100001111;
      square_table[138] = 25'b0111000001001100001101110;
      square_table[139] = 25'b0111000000110001111011111;
      square_table[140] = 25'b0111000000010111101100100;
      square_table[141] = 25'b0110111111111101011111010;
      square_table[142] = 25'b0110111111100011010100011;
      square_table[143] = 25'b0110111111001001001011101;
      square_table[144] = 25'b0110111110101111000101011;
      square_table[145] = 25'b0110111110010101000001011;
      square_table[146] = 25'b0110111101111010111111101;
      square_table[147] = 25'b0110111101100001000000001;
      square_table[148] = 25'b0110111101000111000010111;
      square_table[149] = 25'b0110111100101101001000001;
      square_table[150] = 25'b0110111100010011001111011;
      square_table[151] = 25'b0110111011111001011000111;
      square_table[152] = 25'b0110111011011111100100110;
      square_table[153] = 25'b0110111011000101110010110;
      square_table[154] = 25'b0110111010101100000011001;
      square_table[155] = 25'b0110111010010010010101110;
      square_table[156] = 25'b0110111001111000101010101;
      square_table[157] = 25'b0110111001011111000001101;
      square_table[158] = 25'b0110111001000101011011001;
      square_table[159] = 25'b0110111000101011110110011;
      square_table[160] = 25'b0110111000010010010100010;
      square_table[161] = 25'b0110110111111000110100001;
      square_table[162] = 25'b0110110111011111010110010;
      square_table[163] = 25'b0110110111000101111010111;
      square_table[164] = 25'b0110110110101100100001010;
      square_table[165] = 25'b0110110110010011001010000;
      square_table[166] = 25'b0110110101111001110101001;
      square_table[167] = 25'b0110110101100000100010001;
      square_table[168] = 25'b0110110101000111010001100;
      square_table[169] = 25'b0110110100101110000011010;
      square_table[170] = 25'b0110110100010100110110111;
      square_table[171] = 25'b0110110011111011101100110;
      square_table[172] = 25'b0110110011100010100101000;
      square_table[173] = 25'b0110110011001001011111001;
      square_table[174] = 25'b0110110010110000011011101;
      square_table[175] = 25'b0110110010010111011010010;
      square_table[176] = 25'b0110110001111110011011000;
      square_table[177] = 25'b0110110001100101011110000;
      square_table[178] = 25'b0110110001001100100010111;
      square_table[179] = 25'b0110110000110011101010001;
      square_table[180] = 25'b0110110000011010110011011;
      square_table[181] = 25'b0110110000000001111111000;
      square_table[182] = 25'b0110101111101001001100110;
      square_table[183] = 25'b0110101111010000011100010;
      square_table[184] = 25'b0110101110110111101110010;
      square_table[185] = 25'b0110101110011111000010001;
      square_table[186] = 25'b0110101110000110011000100;
      square_table[187] = 25'b0110101101101101110000101;
      square_table[188] = 25'b0110101101010101001011000;
      square_table[189] = 25'b0110101100111100100111101;
      square_table[190] = 25'b0110101100100100000110001;
      square_table[191] = 25'b0110101100001011100110111;
      square_table[192] = 25'b0110101011110011001001101;
      square_table[193] = 25'b0110101011011010101110011;
      square_table[194] = 25'b0110101011000010010101010;
      square_table[195] = 25'b0110101010101001111110100;
      square_table[196] = 25'b0110101010010001101001100;
      square_table[197] = 25'b0110101001111001010110110;
      square_table[198] = 25'b0110101001100001000110001;
      square_table[199] = 25'b0110101001001000110111010;
      square_table[200] = 25'b0110101000110000101010110;
      square_table[201] = 25'b0110101000011000100000010;
      square_table[202] = 25'b0110101000000000010111111;
      square_table[203] = 25'b0110100111101000010001100;
      square_table[204] = 25'b0110100111010000001101010;
      square_table[205] = 25'b0110100110111000001010111;
      square_table[206] = 25'b0110100110100000001010110;
      square_table[207] = 25'b0110100110001000001100100;
      square_table[208] = 25'b0110100101110000010000011;
      square_table[209] = 25'b0110100101011000010110010;
      square_table[210] = 25'b0110100101000000011110010;
      square_table[211] = 25'b0110100100101000101000000;
      square_table[212] = 25'b0110100100010000110100000;
      square_table[213] = 25'b0110100011111001000010000;
      square_table[214] = 25'b0110100011100001010010001;
      square_table[215] = 25'b0110100011001001100100000;
      square_table[216] = 25'b0110100010110001111000001;
      square_table[217] = 25'b0110100010011010001110000;
      square_table[218] = 25'b0110100010000010100110001;
      square_table[219] = 25'b0110100001101011000000001;
      square_table[220] = 25'b0110100001010011011100001;
      square_table[221] = 25'b0110100000111011111010001;
      square_table[222] = 25'b0110100000100100011010001;
      square_table[223] = 25'b0110100000001100111100010;
      square_table[224] = 25'b0110011111110101100000010;
      square_table[225] = 25'b0110011111011110000110001;
      square_table[226] = 25'b0110011111000110101110010;
      square_table[227] = 25'b0110011110101111011000000;
      square_table[228] = 25'b0110011110011000000011111;
      square_table[229] = 25'b0110011110000000110001110;
      square_table[230] = 25'b0110011101101001100001101;
      square_table[231] = 25'b0110011101010010010011011;
      square_table[232] = 25'b0110011100111011000111010;
      square_table[233] = 25'b0110011100100011111100111;
      square_table[234] = 25'b0110011100001100110100100;
      square_table[235] = 25'b0110011011110101101101111;
      square_table[236] = 25'b0110011011011110101001100;
      square_table[237] = 25'b0110011011000111100110111;
      square_table[238] = 25'b0110011010110000100110010;
      square_table[239] = 25'b0110011010011001100111101;
      square_table[240] = 25'b0110011010000010101010110;
      square_table[241] = 25'b0110011001101011101111111;
      square_table[242] = 25'b0110011001010100110111000;
      square_table[243] = 25'b0110011000111110000000001;
      square_table[244] = 25'b0110011000100111001010111;
      square_table[245] = 25'b0110011000010000010111110;
      square_table[246] = 25'b0110010111111001100110100;
      square_table[247] = 25'b0110010111100010110111001;
      square_table[248] = 25'b0110010111001100001001110;
      square_table[249] = 25'b0110010110110101011110000;
      square_table[250] = 25'b0110010110011110110100100;
      square_table[251] = 25'b0110010110001000001100110;
      square_table[252] = 25'b0110010101110001100110111;
      square_table[253] = 25'b0110010101011011000010110;
      square_table[254] = 25'b0110010101000100100000101;
      square_table[255] = 25'b0110010100101110000000011;
      square_table[256] = 25'b0110010100010111100010000;
      square_table[257] = 25'b0110010100000001000101100;
      square_table[258] = 25'b0110010011101010101011000;
      square_table[259] = 25'b0110010011010100010010001;
      square_table[260] = 25'b0110010010111101111011010;
      square_table[261] = 25'b0110010010100111100110010;
      square_table[262] = 25'b0110010010010001010011000;
      square_table[263] = 25'b0110010001111011000001101;
      square_table[264] = 25'b0110010001100100110010001;
      square_table[265] = 25'b0110010001001110100100100;
      square_table[266] = 25'b0110010000111000011000101;
      square_table[267] = 25'b0110010000100010001110110;
      square_table[268] = 25'b0110010000001100000110101;
      square_table[269] = 25'b0110001111110110000000011;
      square_table[270] = 25'b0110001111011111111011111;
      square_table[271] = 25'b0110001111001001111001010;
      square_table[272] = 25'b0110001110110011111000011;
      square_table[273] = 25'b0110001110011101111001011;
      square_table[274] = 25'b0110001110000111111100001;
      square_table[275] = 25'b0110001101110010000000111;
      square_table[276] = 25'b0110001101011100000111010;
      square_table[277] = 25'b0110001101000110001111100;
      square_table[278] = 25'b0110001100110000011001100;
      square_table[279] = 25'b0110001100011010100101010;
      square_table[280] = 25'b0110001100000100110011001;
      square_table[281] = 25'b0110001011101111000010100;
      square_table[282] = 25'b0110001011011001010011110;
      square_table[283] = 25'b0110001011000011100110101;
      square_table[284] = 25'b0110001010101101111011100;
      square_table[285] = 25'b0110001010011000010010000;
      square_table[286] = 25'b0110001010000010101010100;
      square_table[287] = 25'b0110001001101101000100101;
      square_table[288] = 25'b0110001001010111100000100;
      square_table[289] = 25'b0110001001000001111110010;
      square_table[290] = 25'b0110001000101100011101111;
      square_table[291] = 25'b0110001000010110111111000;
      square_table[292] = 25'b0110001000000001100010000;
      square_table[293] = 25'b0110000111101100000110110;
      square_table[294] = 25'b0110000111010110101101010;
      square_table[295] = 25'b0110000111000001010101100;
      square_table[296] = 25'b0110000110101011111111100;
      square_table[297] = 25'b0110000110010110101011010;
      square_table[298] = 25'b0110000110000001011000110;
      square_table[299] = 25'b0110000101101100001000000;
      square_table[300] = 25'b0110000101010110111001000;
      square_table[301] = 25'b0110000101000001101011110;
      square_table[302] = 25'b0110000100101100100000001;
      square_table[303] = 25'b0110000100010111010110100;
      square_table[304] = 25'b0110000100000010001110010;
      square_table[305] = 25'b0110000011101101000111110;
      square_table[306] = 25'b0110000011011000000011010;
      square_table[307] = 25'b0110000011000011000000010;
      square_table[308] = 25'b0110000010101101111111000;
      square_table[309] = 25'b0110000010011000111111100;
      square_table[310] = 25'b0110000010000100000001111;
      square_table[311] = 25'b0110000001101111000101101;
      square_table[312] = 25'b0110000001011010001011010;
      square_table[313] = 25'b0110000001000101010010100;
      square_table[314] = 25'b0110000000110000011011101;
      square_table[315] = 25'b0110000000011011100110010;
      square_table[316] = 25'b0110000000000110110010110;
      square_table[317] = 25'b0101111111110010000000111;
      square_table[318] = 25'b0101111111011101010000100;
      square_table[319] = 25'b0101111111001000100010000;
      square_table[320] = 25'b0101111110110011110101010;
      square_table[321] = 25'b0101111110011111001001111;
      square_table[322] = 25'b0101111110001010100000011;
      square_table[323] = 25'b0101111101110101111000100;
      square_table[324] = 25'b0101111101100001010010011;
      square_table[325] = 25'b0101111101001100101101110;
      square_table[326] = 25'b0101111100111000001011000;
      square_table[327] = 25'b0101111100100011101001110;
      square_table[328] = 25'b0101111100001111001010010;
      square_table[329] = 25'b0101111011111010101100011;
      square_table[330] = 25'b0101111011100110010000000;
      square_table[331] = 25'b0101111011010001110101011;
      square_table[332] = 25'b0101111010111101011100110;
      square_table[333] = 25'b0101111010101001000101011;
      square_table[334] = 25'b0101111010010100101111101;
      square_table[335] = 25'b0101111010000000011011101;
      square_table[336] = 25'b0101111001101100001001010;
      square_table[337] = 25'b0101111001010111111000100;
      square_table[338] = 25'b0101111001000011101001011;
      square_table[339] = 25'b0101111000101111011011111;
      square_table[340] = 25'b0101111000011011010000000;
      square_table[341] = 25'b0101111000000111000101111;
      square_table[342] = 25'b0101110111110010111101010;
      square_table[343] = 25'b0101110111011110110110001;
      square_table[344] = 25'b0101110111001010110000110;
      square_table[345] = 25'b0101110110110110101101000;
      square_table[346] = 25'b0101110110100010101010111;
      square_table[347] = 25'b0101110110001110101010011;
      square_table[348] = 25'b0101110101111010101011001;
      square_table[349] = 25'b0101110101100110101101111;
      square_table[350] = 25'b0101110101010010110010001;
      square_table[351] = 25'b0101110100111110111000000;
      square_table[352] = 25'b0101110100101010111111100;
      square_table[353] = 25'b0101110100010111001000011;
      square_table[354] = 25'b0101110100000011010011000;
      square_table[355] = 25'b0101110011101111011111010;
      square_table[356] = 25'b0101110011011011101100111;
      square_table[357] = 25'b0101110011000111111100010;
      square_table[358] = 25'b0101110010110100001101001;
      square_table[359] = 25'b0101110010100000011111110;
      square_table[360] = 25'b0101110010001100110011110;
      square_table[361] = 25'b0101110001111001001001010;
      square_table[362] = 25'b0101110001100101100000101;
      square_table[363] = 25'b0101110001010001111001011;
      square_table[364] = 25'b0101110000111110010011110;
      square_table[365] = 25'b0101110000101010101111011;
      square_table[366] = 25'b0101110000010111001100111;
      square_table[367] = 25'b0101110000000011101011111;
      square_table[368] = 25'b0101101111110000001100011;
      square_table[369] = 25'b0101101111011100101110101;
      square_table[370] = 25'b0101101111001001010010001;
      square_table[371] = 25'b0101101110110101110111010;
      square_table[372] = 25'b0101101110100010011110000;
      square_table[373] = 25'b0101101110001111000110010;
      square_table[374] = 25'b0101101101111011110000001;
      square_table[375] = 25'b0101101101101000011011011;
      square_table[376] = 25'b0101101101010101001000001;
      square_table[377] = 25'b0101101101000001110110100;
      square_table[378] = 25'b0101101100101110100110011;
      square_table[379] = 25'b0101101100011011010111111;
      square_table[380] = 25'b0101101100001000001010111;
      square_table[381] = 25'b0101101011110100111111010;
      square_table[382] = 25'b0101101011100001110101010;
      square_table[383] = 25'b0101101011001110101100110;
      square_table[384] = 25'b0101101010111011100101110;
      square_table[385] = 25'b0101101010101000100000001;
      square_table[386] = 25'b0101101010010101011100011;
      square_table[387] = 25'b0101101010000010011001111;
      square_table[388] = 25'b0101101001101111011000101;
      square_table[389] = 25'b0101101001011100011001010;
      square_table[390] = 25'b0101101001001001011011010;
      square_table[391] = 25'b0101101000110110011110110;
      square_table[392] = 25'b0101101000100011100011110;
      square_table[393] = 25'b0101101000010000101010001;
      square_table[394] = 25'b0101100111111101110010010;
      square_table[395] = 25'b0101100111101010111011110;
      square_table[396] = 25'b0101100111011000000110100;
      square_table[397] = 25'b0101100111000101010010110;
      square_table[398] = 25'b0101100110110010100000111;
      square_table[399] = 25'b0101100110011111110000001;
      square_table[400] = 25'b0101100110001101000001000;
      square_table[401] = 25'b0101100101111010010011010;
      square_table[402] = 25'b0101100101100111100110111;
      square_table[403] = 25'b0101100101010100111100010;
      square_table[404] = 25'b0101100101000010010010111;
      square_table[405] = 25'b0101100100101111101011000;
      square_table[406] = 25'b0101100100011101000100100;
      square_table[407] = 25'b0101100100001010011111101;
      square_table[408] = 25'b0101100011110111111100001;
      square_table[409] = 25'b0101100011100101011010000;
      square_table[410] = 25'b0101100011010010111001011;
      square_table[411] = 25'b0101100011000000011010011;
      square_table[412] = 25'b0101100010101101111100101;
      square_table[413] = 25'b0101100010011011100000011;
      square_table[414] = 25'b0101100010001001000101011;
      square_table[415] = 25'b0101100001110110101100000;
      square_table[416] = 25'b0101100001100100010100001;
      square_table[417] = 25'b0101100001010001111101100;
      square_table[418] = 25'b0101100000111111101000100;
      square_table[419] = 25'b0101100000101101010100101;
      square_table[420] = 25'b0101100000011011000010011;
      square_table[421] = 25'b0101100000001000110001101;
      square_table[422] = 25'b0101011111110110100010010;
      square_table[423] = 25'b0101011111100100010100010;
      square_table[424] = 25'b0101011111010010000111101;
      square_table[425] = 25'b0101011110111111111100011;
      square_table[426] = 25'b0101011110101101110010110;
      square_table[427] = 25'b0101011110011011101010011;
      square_table[428] = 25'b0101011110001001100011011;
      square_table[429] = 25'b0101011101110111011101111;
      square_table[430] = 25'b0101011101100101011001101;
      square_table[431] = 25'b0101011101010011010110111;
      square_table[432] = 25'b0101011101000001010101011;
      square_table[433] = 25'b0101011100101111010101100;
      square_table[434] = 25'b0101011100011101010111000;
      square_table[435] = 25'b0101011100001011011001111;
      square_table[436] = 25'b0101011011111001011110000;
      square_table[437] = 25'b0101011011100111100011101;
      square_table[438] = 25'b0101011011010101101010100;
      square_table[439] = 25'b0101011011000011110010111;
      square_table[440] = 25'b0101011010110001111100100;
      square_table[441] = 25'b0101011010100000000111110;
      square_table[442] = 25'b0101011010001110010100001;
      square_table[443] = 25'b0101011001111100100010000;
      square_table[444] = 25'b0101011001101010110001010;
      square_table[445] = 25'b0101011001011001000010000;
      square_table[446] = 25'b0101011001000111010011111;
      square_table[447] = 25'b0101011000110101100111001;
      square_table[448] = 25'b0101011000100011111011111;
      square_table[449] = 25'b0101011000010010010001111;
      square_table[450] = 25'b0101011000000000101001011;
      square_table[451] = 25'b0101010111101111000010001;
      square_table[452] = 25'b0101010111011101011100001;
      square_table[453] = 25'b0101010111001011110111100;
      square_table[454] = 25'b0101010110111010010100011;
      square_table[455] = 25'b0101010110101000110010100;
      square_table[456] = 25'b0101010110010111010010000;
      square_table[457] = 25'b0101010110000101110010110;
      square_table[458] = 25'b0101010101110100010101000;
      square_table[459] = 25'b0101010101100010111000100;
      square_table[460] = 25'b0101010101010001011101010;
      square_table[461] = 25'b0101010101000000000011100;
      square_table[462] = 25'b0101010100101110101010111;
      square_table[463] = 25'b0101010100011101010011111;
      square_table[464] = 25'b0101010100001011111110000;
      square_table[465] = 25'b0101010011111010101001100;
      square_table[466] = 25'b0101010011101001010110010;
      square_table[467] = 25'b0101010011011000000100011;
      square_table[468] = 25'b0101010011000110110011110;
      square_table[469] = 25'b0101010010110101100100101;
      square_table[470] = 25'b0101010010100100010110110;
      square_table[471] = 25'b0101010010010011001010001;
      square_table[472] = 25'b0101010010000001111110110;
      square_table[473] = 25'b0101010001110000110100111;
      square_table[474] = 25'b0101010001011111101100001;
      square_table[475] = 25'b0101010001001110100100110;
      square_table[476] = 25'b0101010000111101011110100;
      square_table[477] = 25'b0101010000101100011001110;
      square_table[478] = 25'b0101010000011011010110010;
      square_table[479] = 25'b0101010000001010010100000;
      square_table[480] = 25'b0101001111111001010011010;
      square_table[481] = 25'b0101001111101000010011101;
      square_table[482] = 25'b0101001111010111010101011;
      square_table[483] = 25'b0101001111000110011000010;
      square_table[484] = 25'b0101001110110101011100101;
      square_table[485] = 25'b0101001110100100100010000;
      square_table[486] = 25'b0101001110010011101000110;
      square_table[487] = 25'b0101001110000010110001000;
      square_table[488] = 25'b0101001101110001111010011;
      square_table[489] = 25'b0101001101100001000101000;
      square_table[490] = 25'b0101001101010000010000110;
      square_table[491] = 25'b0101001100111111011110000;
      square_table[492] = 25'b0101001100101110101100101;
      square_table[493] = 25'b0101001100011101111100010;
      square_table[494] = 25'b0101001100001101001101010;
      square_table[495] = 25'b0101001011111100011111101;
      square_table[496] = 25'b0101001011101011110010111;
      square_table[497] = 25'b0101001011011011000111111;
      square_table[498] = 25'b0101001011001010011101111;
      square_table[499] = 25'b0101001010111001110101000;
      square_table[500] = 25'b0101001010101001001101101;
      square_table[501] = 25'b0101001010011000100111100;
      square_table[502] = 25'b0101001010001000000010100;
      square_table[503] = 25'b0101001001110111011110111;
      square_table[504] = 25'b0101001001100110111100010;
      square_table[505] = 25'b0101001001010110011011000;
      square_table[506] = 25'b0101001001000101111011001;
      square_table[507] = 25'b0101001000110101011100010;
      square_table[508] = 25'b0101001000100100111110111;
      square_table[509] = 25'b0101001000010100100010101;
      square_table[510] = 25'b0101001000000100000111101;
      square_table[511] = 25'b0101000111110011101101110;
      square_table[512] = 25'b0101000111100011010101001;
      square_table[513] = 25'b0101000111010010111101110;
      square_table[514] = 25'b0101000111000010100111101;
      square_table[515] = 25'b0101000110110010010010111;
      square_table[516] = 25'b0101000110100001111111000;
      square_table[517] = 25'b0101000110010001101100110;
      square_table[518] = 25'b0101000110000001011011011;
      square_table[519] = 25'b0101000101110001001011011;
      square_table[520] = 25'b0101000101100000111100101;
      square_table[521] = 25'b0101000101010000101111001;
      square_table[522] = 25'b0101000101000000100010100;
      square_table[523] = 25'b0101000100110000010111011;
      square_table[524] = 25'b0101000100100000001101011;
      square_table[525] = 25'b0101000100010000000100101;
      square_table[526] = 25'b0101000011111111111101001;
      square_table[527] = 25'b0101000011101111110110110;
      square_table[528] = 25'b0101000011011111110001101;
      square_table[529] = 25'b0101000011001111101101101;
      square_table[530] = 25'b0101000010111111101010110;
      square_table[531] = 25'b0101000010101111101001011;
      square_table[532] = 25'b0101000010011111101001000;
      square_table[533] = 25'b0101000010001111101001111;
      square_table[534] = 25'b0101000001111111101011110;
      square_table[535] = 25'b0101000001101111101111000;
      square_table[536] = 25'b0101000001011111110011011;
      square_table[537] = 25'b0101000001001111111000111;
      square_table[538] = 25'b0101000000111111111111101;
      square_table[539] = 25'b0101000000110000000111100;
      square_table[540] = 25'b0101000000100000010000101;
      square_table[541] = 25'b0101000000010000011010111;
      square_table[542] = 25'b0101000000000000100110011;
      square_table[543] = 25'b0100111111110000110011000;
      square_table[544] = 25'b0100111111100001000000101;
      square_table[545] = 25'b0100111111010001001111101;
      square_table[546] = 25'b0100111111000001011111111;
      square_table[547] = 25'b0100111110110001110001000;
      square_table[548] = 25'b0100111110100010000011100;
      square_table[549] = 25'b0100111110010010010111001;
      square_table[550] = 25'b0100111110000010101100000;
      square_table[551] = 25'b0100111101110011000001111;
      square_table[552] = 25'b0100111101100011011000111;
      square_table[553] = 25'b0100111101010011110001001;
      square_table[554] = 25'b0100111101000100001010100;
      square_table[555] = 25'b0100111100110100100101000;
      square_table[556] = 25'b0100111100100101000000110;
      square_table[557] = 25'b0100111100010101011101101;
      square_table[558] = 25'b0100111100000101111011100;
      square_table[559] = 25'b0100111011110110011010110;
      square_table[560] = 25'b0100111011100110111010111;
      square_table[561] = 25'b0100111011010111011100010;
      square_table[562] = 25'b0100111011000111111110110;
      square_table[563] = 25'b0100111010111000100010100;
      square_table[564] = 25'b0100111010101001000111011;
      square_table[565] = 25'b0100111010011001101101011;
      square_table[566] = 25'b0100111010001010010100011;
      square_table[567] = 25'b0100111001111010111100100;
      square_table[568] = 25'b0100111001101011100110000;
      square_table[569] = 25'b0100111001011100010000011;
      square_table[570] = 25'b0100111001001100111100000;
      square_table[571] = 25'b0100111000111101101000101;
      square_table[572] = 25'b0100111000101110010110100;
      square_table[573] = 25'b0100111000011111000101011;
      square_table[574] = 25'b0100111000001111110101100;
      square_table[575] = 25'b0100111000000000100110101;
      square_table[576] = 25'b0100110111110001011001000;
      square_table[577] = 25'b0100110111100010001100010;
      square_table[578] = 25'b0100110111010011000000111;
      square_table[579] = 25'b0100110111000011110110100;
      square_table[580] = 25'b0100110110110100101101010;
      square_table[581] = 25'b0100110110100101100101001;
      square_table[582] = 25'b0100110110010110011110000;
      square_table[583] = 25'b0100110110000111011000000;
      square_table[584] = 25'b0100110101111000010011001;
      square_table[585] = 25'b0100110101101001001111011;
      square_table[586] = 25'b0100110101011010001100111;
      square_table[587] = 25'b0100110101001011001011010;
      square_table[588] = 25'b0100110100111100001010110;
      square_table[589] = 25'b0100110100101101001011011;
      square_table[590] = 25'b0100110100011110001101001;
      square_table[591] = 25'b0100110100001111001111111;
      square_table[592] = 25'b0100110100000000010011110;
      square_table[593] = 25'b0100110011110001011000110;
      square_table[594] = 25'b0100110011100010011110110;
      square_table[595] = 25'b0100110011010011100101111;
      square_table[596] = 25'b0100110011000100101110001;
      square_table[597] = 25'b0100110010110101110111100;
      square_table[598] = 25'b0100110010100111000001110;
      square_table[599] = 25'b0100110010011000001101011;
      square_table[600] = 25'b0100110010001001011001110;
      square_table[601] = 25'b0100110001111010100111100;
      square_table[602] = 25'b0100110001101011110110001;
      square_table[603] = 25'b0100110001011101000101111;
      square_table[604] = 25'b0100110001001110010110110;
      square_table[605] = 25'b0100110000111111101000101;
      square_table[606] = 25'b0100110000110000111011100;
      square_table[607] = 25'b0100110000100010001111011;
      square_table[608] = 25'b0100110000010011100100101;
      square_table[609] = 25'b0100110000000100111010110;
      square_table[610] = 25'b0100101111110110010001111;
      square_table[611] = 25'b0100101111100111101010000;
      square_table[612] = 25'b0100101111011001000011011;
      square_table[613] = 25'b0100101111001010011101110;
      square_table[614] = 25'b0100101110111011111001001;
      square_table[615] = 25'b0100101110101101010101101;
      square_table[616] = 25'b0100101110011110110011000;
      square_table[617] = 25'b0100101110010000010001100;
      square_table[618] = 25'b0100101110000001110001001;
      square_table[619] = 25'b0100101101110011010001111;
      square_table[620] = 25'b0100101101100100110011101;
      square_table[621] = 25'b0100101101010110010110010;
      square_table[622] = 25'b0100101101000111111001111;
      square_table[623] = 25'b0100101100111001011110110;
      square_table[624] = 25'b0100101100101011000100110;
      square_table[625] = 25'b0100101100011100101011100;
      square_table[626] = 25'b0100101100001110010011011;
      square_table[627] = 25'b0100101011111111111100011;
      square_table[628] = 25'b0100101011110001100110010;
      square_table[629] = 25'b0100101011100011010001011;
      square_table[630] = 25'b0100101011010100111101011;
      square_table[631] = 25'b0100101011000110101010010;
      square_table[632] = 25'b0100101010111000011000011;
      square_table[633] = 25'b0100101010101010000111100;
      square_table[634] = 25'b0100101010011011110111100;
      square_table[635] = 25'b0100101010001101101000101;
      square_table[636] = 25'b0100101001111111011011000;
      square_table[637] = 25'b0100101001110001001101111;
      square_table[638] = 25'b0100101001100011000010010;
      square_table[639] = 25'b0100101001010100110111011;
      square_table[640] = 25'b0100101001000110101101100;
      square_table[641] = 25'b0100101000111000100100111;
      square_table[642] = 25'b0100101000101010011101000;
      square_table[643] = 25'b0100101000011100010110001;
      square_table[644] = 25'b0100101000001110010000100;
      square_table[645] = 25'b0100101000000000001011101;
      square_table[646] = 25'b0100100111110010001000000;
      square_table[647] = 25'b0100100111100100000101001;
      square_table[648] = 25'b0100100111010110000011100;
      square_table[649] = 25'b0100100111001000000010101;
      square_table[650] = 25'b0100100110111010000010111;
      square_table[651] = 25'b0100100110101100000100001;
      square_table[652] = 25'b0100100110011110000110011;
      square_table[653] = 25'b0100100110010000001001101;
      square_table[654] = 25'b0100100110000010001101111;
      square_table[655] = 25'b0100100101110100010011000;
      square_table[656] = 25'b0100100101100110011001010;
      square_table[657] = 25'b0100100101011000100000011;
      square_table[658] = 25'b0100100101001010101000011;
      square_table[659] = 25'b0100100100111100110001100;
      square_table[660] = 25'b0100100100101110111011110;
      square_table[661] = 25'b0100100100100001000110111;
      square_table[662] = 25'b0100100100010011010010111;
      square_table[663] = 25'b0100100100000101100000000;
      square_table[664] = 25'b0100100011110111101110001;
      square_table[665] = 25'b0100100011101001111101000;
      square_table[666] = 25'b0100100011011100001101001;
      square_table[667] = 25'b0100100011001110011101111;
      square_table[668] = 25'b0100100011000000101111111;
      square_table[669] = 25'b0100100010110011000010111;
      square_table[670] = 25'b0100100010100101010110110;
      square_table[671] = 25'b0100100010010111101011100;
      square_table[672] = 25'b0100100010001010000001010;
      square_table[673] = 25'b0100100001111100011000000;
      square_table[674] = 25'b0100100001101110101111110;
      square_table[675] = 25'b0100100001100001001000100;
      square_table[676] = 25'b0100100001010011100010000;
      square_table[677] = 25'b0100100001000101111100101;
      square_table[678] = 25'b0100100000111000011000010;
      square_table[679] = 25'b0100100000101010110100110;
      square_table[680] = 25'b0100100000011101010010010;
      square_table[681] = 25'b0100100000001111110000101;
      square_table[682] = 25'b0100100000000010010000000;
      square_table[683] = 25'b0100011111110100110000010;
      square_table[684] = 25'b0100011111100111010001101;
      square_table[685] = 25'b0100011111011001110011111;
      square_table[686] = 25'b0100011111001100010111000;
      square_table[687] = 25'b0100011110111110111011000;
      square_table[688] = 25'b0100011110110001100000000;
      square_table[689] = 25'b0100011110100100000110001;
      square_table[690] = 25'b0100011110010110101101000;
      square_table[691] = 25'b0100011110001001010100111;
      square_table[692] = 25'b0100011101111011111101110;
      square_table[693] = 25'b0100011101101110100111011;
      square_table[694] = 25'b0100011101100001010010000;
      square_table[695] = 25'b0100011101010011111101110;
      square_table[696] = 25'b0100011101000110101010001;
      square_table[697] = 25'b0100011100111001010111101;
      square_table[698] = 25'b0100011100101100000110001;
      square_table[699] = 25'b0100011100011110110101011;
      square_table[700] = 25'b0100011100010001100101101;
      square_table[701] = 25'b0100011100000100010110110;
      square_table[702] = 25'b0100011011110111001000111;
      square_table[703] = 25'b0100011011101001111100000;
      square_table[704] = 25'b0100011011011100101111111;
      square_table[705] = 25'b0100011011001111100100110;
      square_table[706] = 25'b0100011011000010011010100;
      square_table[707] = 25'b0100011010110101010001001;
      square_table[708] = 25'b0100011010101000001000111;
      square_table[709] = 25'b0100011010011011000001010;
      square_table[710] = 25'b0100011010001101111010110;
      square_table[711] = 25'b0100011010000000110101000;
      square_table[712] = 25'b0100011001110011110000011;
      square_table[713] = 25'b0100011001100110101100100;
      square_table[714] = 25'b0100011001011001101001100;
      square_table[715] = 25'b0100011001001100100111101;
      square_table[716] = 25'b0100011000111111100110100;
      square_table[717] = 25'b0100011000110010100110010;
      square_table[718] = 25'b0100011000100101100111000;
      square_table[719] = 25'b0100011000011000101000100;
      square_table[720] = 25'b0100011000001011101010111;
      square_table[721] = 25'b0100010111111110101110011;
      square_table[722] = 25'b0100010111110001110010101;
      square_table[723] = 25'b0100010111100100110111111;
      square_table[724] = 25'b0100010111010111111110000;
      square_table[725] = 25'b0100010111001011000100111;
      square_table[726] = 25'b0100010110111110001100110;
      square_table[727] = 25'b0100010110110001010101100;
      square_table[728] = 25'b0100010110100100011111001;
      square_table[729] = 25'b0100010110010111101001110;
      square_table[730] = 25'b0100010110001010110101001;
      square_table[731] = 25'b0100010101111110000001011;
      square_table[732] = 25'b0100010101110001001110101;
      square_table[733] = 25'b0100010101100100011100101;
      square_table[734] = 25'b0100010101010111101011100;
      square_table[735] = 25'b0100010101001010111011011;
      square_table[736] = 25'b0100010100111110001100001;
      square_table[737] = 25'b0100010100110001011101110;
      square_table[738] = 25'b0100010100100100110000001;
      square_table[739] = 25'b0100010100011000000011101;
      square_table[740] = 25'b0100010100001011010111110;
      square_table[741] = 25'b0100010011111110101100111;
      square_table[742] = 25'b0100010011110010000010111;
      square_table[743] = 25'b0100010011100101011001101;
      square_table[744] = 25'b0100010011011000110001011;
      square_table[745] = 25'b0100010011001100001001110;
      square_table[746] = 25'b0100010010111111100011011;
      square_table[747] = 25'b0100010010110010111101101;
      square_table[748] = 25'b0100010010100110011000110;
      square_table[749] = 25'b0100010010011001110100110;
      square_table[750] = 25'b0100010010001101010001110;
      square_table[751] = 25'b0100010010000000101111100;
      square_table[752] = 25'b0100010001110100001110000;
      square_table[753] = 25'b0100010001100111101101101;
      square_table[754] = 25'b0100010001011011001101110;
      square_table[755] = 25'b0100010001001110101111000;
      square_table[756] = 25'b0100010001000010010001000;
      square_table[757] = 25'b0100010000110101110011111;
      square_table[758] = 25'b0100010000101001010111101;
      square_table[759] = 25'b0100010000011100111100010;
      square_table[760] = 25'b0100010000010000100001110;
      square_table[761] = 25'b0100010000000100001000000;
      square_table[762] = 25'b0100001111110111101111010;
      square_table[763] = 25'b0100001111101011010111000;
      square_table[764] = 25'b0100001111011110111111111;
      square_table[765] = 25'b0100001111010010101001101;
      square_table[766] = 25'b0100001111000110010100001;
      square_table[767] = 25'b0100001110111001111111100;
      square_table[768] = 25'b0100001110101101101011110;
      square_table[769] = 25'b0100001110100001011000110;
      square_table[770] = 25'b0100001110010101000110100;
      square_table[771] = 25'b0100001110001000110101010;
      square_table[772] = 25'b0100001101111100100100101;
      square_table[773] = 25'b0100001101110000010101001;
      square_table[774] = 25'b0100001101100100000110010;
      square_table[775] = 25'b0100001101010111111000011;
      square_table[776] = 25'b0100001101001011101011001;
      square_table[777] = 25'b0100001100111111011110111;
      square_table[778] = 25'b0100001100110011010011100;
      square_table[779] = 25'b0100001100100111001000110;
      square_table[780] = 25'b0100001100011010111111000;
      square_table[781] = 25'b0100001100001110110110000;
      square_table[782] = 25'b0100001100000010101101111;
      square_table[783] = 25'b0100001011110110100110011;
      square_table[784] = 25'b0100001011101010011111111;
      square_table[785] = 25'b0100001011011110011010001;
      square_table[786] = 25'b0100001011010010010101010;
      square_table[787] = 25'b0100001011000110010001010;
      square_table[788] = 25'b0100001010111010001110000;
      square_table[789] = 25'b0100001010101110001011100;
      square_table[790] = 25'b0100001010100010001001111;
      square_table[791] = 25'b0100001010010110001001001;
      square_table[792] = 25'b0100001010001010001001001;
      square_table[793] = 25'b0100001001111110001001111;
      square_table[794] = 25'b0100001001110010001011100;
      square_table[795] = 25'b0100001001100110001110000;
      square_table[796] = 25'b0100001001011010010001010;
      square_table[797] = 25'b0100001001001110010101010;
      square_table[798] = 25'b0100001001000010011001111;
      square_table[799] = 25'b0100001000110110011111101;
      square_table[800] = 25'b0100001000101010100110001;
      square_table[801] = 25'b0100001000011110101101011;
      square_table[802] = 25'b0100001000010010110101011;
      square_table[803] = 25'b0100001000000110111110011;
      square_table[804] = 25'b0100000111111011000111111;
      square_table[805] = 25'b0100000111101111010010011;
      square_table[806] = 25'b0100000111100011011101101;
      square_table[807] = 25'b0100000111010111101001100;
      square_table[808] = 25'b0100000111001011110110100;
      square_table[809] = 25'b0100000111000000000100000;
      square_table[810] = 25'b0100000110110100010010100;
      square_table[811] = 25'b0100000110101000100001101;
      square_table[812] = 25'b0100000110011100110001110;
      square_table[813] = 25'b0100000110010001000010100;
      square_table[814] = 25'b0100000110000101010100000;
      square_table[815] = 25'b0100000101111001100110011;
      square_table[816] = 25'b0100000101101101111001100;
      square_table[817] = 25'b0100000101100010001101011;
      square_table[818] = 25'b0100000101010110100010001;
      square_table[819] = 25'b0100000101001010110111101;
      square_table[820] = 25'b0100000100111111001110000;
      square_table[821] = 25'b0100000100110011100100111;
      square_table[822] = 25'b0100000100100111111100110;
      square_table[823] = 25'b0100000100011100010101011;
      square_table[824] = 25'b0100000100010000101110110;
      square_table[825] = 25'b0100000100000101001000111;
      square_table[826] = 25'b0100000011111001100011111;
      square_table[827] = 25'b0100000011101101111111100;
      square_table[828] = 25'b0100000011100010011100000;
      square_table[829] = 25'b0100000011010110111001010;
      square_table[830] = 25'b0100000011001011010111011;
      square_table[831] = 25'b0100000010111111110110000;
      square_table[832] = 25'b0100000010110100010101101;
      square_table[833] = 25'b0100000010101000110101111;
      square_table[834] = 25'b0100000010011101010111000;
      square_table[835] = 25'b0100000010010001111000110;
      square_table[836] = 25'b0100000010000110011011011;
      square_table[837] = 25'b0100000001111010111110110;
      square_table[838] = 25'b0100000001101111100011000;
      square_table[839] = 25'b0100000001100100000111110;
      square_table[840] = 25'b0100000001011000101101101;
      square_table[841] = 25'b0100000001001101010011111;
      square_table[842] = 25'b0100000001000001111011001;
      square_table[843] = 25'b0100000000110110100011000;
      square_table[844] = 25'b0100000000101011001011110;
      square_table[845] = 25'b0100000000011111110101010;
      square_table[846] = 25'b0100000000010100011111011;
      square_table[847] = 25'b0100000000001001001010010;
      square_table[848] = 25'b0011111111111101110101111;
      square_table[849] = 25'b0011111111110010100010011;
      square_table[850] = 25'b0011111111100111001111100;
      square_table[851] = 25'b0011111111011011111101100;
      square_table[852] = 25'b0011111111010000101100001;
      square_table[853] = 25'b0011111111000101011011100;
      square_table[854] = 25'b0011111110111010001011110;
      square_table[855] = 25'b0011111110101110111100101;
      square_table[856] = 25'b0011111110100011101110011;
      square_table[857] = 25'b0011111110011000100000110;
      square_table[858] = 25'b0011111110001101010100000;
      square_table[859] = 25'b0011111110000010000111111;
      square_table[860] = 25'b0011111101110110111100100;
      square_table[861] = 25'b0011111101101011110001110;
      square_table[862] = 25'b0011111101100000100111111;
      square_table[863] = 25'b0011111101010101011110110;
      square_table[864] = 25'b0011111101001010010110010;
      square_table[865] = 25'b0011111100111111001110101;
      square_table[866] = 25'b0011111100110100000111100;
      square_table[867] = 25'b0011111100101001000001011;
      square_table[868] = 25'b0011111100011101111011111;
      square_table[869] = 25'b0011111100010010110111001;
      square_table[870] = 25'b0011111100000111110011001;
      square_table[871] = 25'b0011111011111100101111110;
      square_table[872] = 25'b0011111011110001101101001;
      square_table[873] = 25'b0011111011100110101011010;
      square_table[874] = 25'b0011111011011011101010001;
      square_table[875] = 25'b0011111011010000101001101;
      square_table[876] = 25'b0011111011000101101001111;
      square_table[877] = 25'b0011111010111010101010111;
      square_table[878] = 25'b0011111010101111101100110;
      square_table[879] = 25'b0011111010100100101111010;
      square_table[880] = 25'b0011111010011001110010011;
      square_table[881] = 25'b0011111010001110110110011;
      square_table[882] = 25'b0011111010000011111010111;
      square_table[883] = 25'b0011111001111001000000010;
      square_table[884] = 25'b0011111001101110000110010;
      square_table[885] = 25'b0011111001100011001101001;
      square_table[886] = 25'b0011111001011000010100100;
      square_table[887] = 25'b0011111001001101011100110;
      square_table[888] = 25'b0011111001000010100101101;
      square_table[889] = 25'b0011111000110111101111001;
      square_table[890] = 25'b0011111000101100111001100;
      square_table[891] = 25'b0011111000100010000100100;
      square_table[892] = 25'b0011111000010111010000010;
      square_table[893] = 25'b0011111000001100011100101;
      square_table[894] = 25'b0011111000000001101001110;
      square_table[895] = 25'b0011110111110110110111101;
      square_table[896] = 25'b0011110111101100000110010;
      square_table[897] = 25'b0011110111100001010101011;
      square_table[898] = 25'b0011110111010110100101011;
      square_table[899] = 25'b0011110111001011110110000;
      square_table[900] = 25'b0011110111000001000111010;
      square_table[901] = 25'b0011110110110110011001011;
      square_table[902] = 25'b0011110110101011101100001;
      square_table[903] = 25'b0011110110100000111111101;
      square_table[904] = 25'b0011110110010110010011110;
      square_table[905] = 25'b0011110110001011101000100;
      square_table[906] = 25'b0011110110000000111110001;
      square_table[907] = 25'b0011110101110110010100010;
      square_table[908] = 25'b0011110101101011101011010;
      square_table[909] = 25'b0011110101100001000010110;
      square_table[910] = 25'b0011110101010110011011000;
      square_table[911] = 25'b0011110101001011110100001;
      square_table[912] = 25'b0011110101000001001101101;
      square_table[913] = 25'b0011110100110110101000000;
      square_table[914] = 25'b0011110100101100000011001;
      square_table[915] = 25'b0011110100100001011110110;
      square_table[916] = 25'b0011110100010110111011010;
      square_table[917] = 25'b0011110100001100011000011;
      square_table[918] = 25'b0011110100000001110110001;
      square_table[919] = 25'b0011110011110111010100101;
      square_table[920] = 25'b0011110011101100110011101;
      square_table[921] = 25'b0011110011100010010011011;
      square_table[922] = 25'b0011110011010111110100000;
      square_table[923] = 25'b0011110011001101010101010;
      square_table[924] = 25'b0011110011000010110111001;
      square_table[925] = 25'b0011110010111000011001100;
      square_table[926] = 25'b0011110010101101111100110;
      square_table[927] = 25'b0011110010100011100000101;
      square_table[928] = 25'b0011110010011001000101010;
      square_table[929] = 25'b0011110010001110101010100;
      square_table[930] = 25'b0011110010000100010000010;
      square_table[931] = 25'b0011110001111001110110110;
      square_table[932] = 25'b0011110001101111011110000;
      square_table[933] = 25'b0011110001100101000110000;
      square_table[934] = 25'b0011110001011010101110101;
      square_table[935] = 25'b0011110001010000010111110;
      square_table[936] = 25'b0011110001000110000001110;
      square_table[937] = 25'b0011110000111011101100001;
      square_table[938] = 25'b0011110000110001010111100;
      square_table[939] = 25'b0011110000100111000011011;
      square_table[940] = 25'b0011110000011100101111111;
      square_table[941] = 25'b0011110000010010011101001;
      square_table[942] = 25'b0011110000001000001011000;
      square_table[943] = 25'b0011101111111101111001100;
      square_table[944] = 25'b0011101111110011101000110;
      square_table[945] = 25'b0011101111101001011000100;
      square_table[946] = 25'b0011101111011111001001000;
      square_table[947] = 25'b0011101111010100111010011;
      square_table[948] = 25'b0011101111001010101100001;
      square_table[949] = 25'b0011101111000000011110100;
      square_table[950] = 25'b0011101110110110010001110;
      square_table[951] = 25'b0011101110101100000101100;
      square_table[952] = 25'b0011101110100001111010000;
      square_table[953] = 25'b0011101110010111101111000;
      square_table[954] = 25'b0011101110001101100100111;
      square_table[955] = 25'b0011101110000011011011010;
      square_table[956] = 25'b0011101101111001010010010;
      square_table[957] = 25'b0011101101101111001001111;
      square_table[958] = 25'b0011101101100101000010001;
      square_table[959] = 25'b0011101101011010111011001;
      square_table[960] = 25'b0011101101010000110100111;
      square_table[961] = 25'b0011101101000110101111001;
      square_table[962] = 25'b0011101100111100101010000;
      square_table[963] = 25'b0011101100110010100101101;
      square_table[964] = 25'b0011101100101000100001101;
      square_table[965] = 25'b0011101100011110011110100;
      square_table[966] = 25'b0011101100010100011100000;
      square_table[967] = 25'b0011101100001010011010001;
      square_table[968] = 25'b0011101100000000011000111;
      square_table[969] = 25'b0011101011110110011000010;
      square_table[970] = 25'b0011101011101100011000011;
      square_table[971] = 25'b0011101011100010011001000;
      square_table[972] = 25'b0011101011011000011010010;
      square_table[973] = 25'b0011101011001110011100010;
      square_table[974] = 25'b0011101011000100011110110;
      square_table[975] = 25'b0011101010111010100001111;
      square_table[976] = 25'b0011101010110000100101110;
      square_table[977] = 25'b0011101010100110101010010;
      square_table[978] = 25'b0011101010011100101111011;
      square_table[979] = 25'b0011101010010010110101001;
      square_table[980] = 25'b0011101010001000111011011;
      square_table[981] = 25'b0011101001111111000010011;
      square_table[982] = 25'b0011101001110101001010000;
      square_table[983] = 25'b0011101001101011010010010;
      square_table[984] = 25'b0011101001100001011011000;
      square_table[985] = 25'b0011101001010111100100100;
      square_table[986] = 25'b0011101001001101101110101;
      square_table[987] = 25'b0011101001000011111001011;
      square_table[988] = 25'b0011101000111010000100101;
      square_table[989] = 25'b0011101000110000010000101;
      square_table[990] = 25'b0011101000100110011101010;
      square_table[991] = 25'b0011101000011100101010100;
      square_table[992] = 25'b0011101000010010111000010;
      square_table[993] = 25'b0011101000001001000110101;
      square_table[994] = 25'b0011100111111111010101110;
      square_table[995] = 25'b0011100111110101100101100;
      square_table[996] = 25'b0011100111101011110101110;
      square_table[997] = 25'b0011100111100010000110101;
      square_table[998] = 25'b0011100111011000011000000;
      square_table[999] = 25'b0011100111001110101010011;
      square_table[1000] = 25'b0011100111000100111101000;
      square_table[1001] = 25'b0011100110111011010000011;
      square_table[1002] = 25'b0011100110110001100100010;
      square_table[1003] = 25'b0011100110100111111000110;
      square_table[1004] = 25'b0011100110011110001110001;
      square_table[1005] = 25'b0011100110010100100011110;
      square_table[1006] = 25'b0011100110001010111010001;
      square_table[1007] = 25'b0011100110000001010001010;
      square_table[1008] = 25'b0011100101110111101000111;
      square_table[1009] = 25'b0011100101101110000001000;
      square_table[1010] = 25'b0011100101100100011001111;
      square_table[1011] = 25'b0011100101011010110011010;
      square_table[1012] = 25'b0011100101010001001101010;
      square_table[1013] = 25'b0011100101000111100111111;
      square_table[1014] = 25'b0011100100111110000011000;
      square_table[1015] = 25'b0011100100110100011110111;
      square_table[1016] = 25'b0011100100101010111011011;
      square_table[1017] = 25'b0011100100100001011000011;
      square_table[1018] = 25'b0011100100010111110101111;
      square_table[1019] = 25'b0011100100001110010100010;
      square_table[1020] = 25'b0011100100000100110011000;
      square_table[1021] = 25'b0011100011111011010010011;
      square_table[1022] = 25'b0011100011110001110010100;
      square_table[1023] = 25'b0011100011101000010011000;
      square_table[1024] = 25'b0011100011011110110100010;
      square_table[1025] = 25'b0011100011010101010110000;
      square_table[1026] = 25'b0011100011001011111000011;
      square_table[1027] = 25'b0011100011000010011011010;
      square_table[1028] = 25'b0011100010111000111110111;
      square_table[1029] = 25'b0011100010101111100011000;
      square_table[1030] = 25'b0011100010100110000111110;
      square_table[1031] = 25'b0011100010011100101101001;
      square_table[1032] = 25'b0011100010010011010011000;
      square_table[1033] = 25'b0011100010001001111001100;
      square_table[1034] = 25'b0011100010000000100000100;
      square_table[1035] = 25'b0011100001110111001000010;
      square_table[1036] = 25'b0011100001101101110000011;
      square_table[1037] = 25'b0011100001100100011001010;
      square_table[1038] = 25'b0011100001011011000010101;
      square_table[1039] = 25'b0011100001010001101100101;
      square_table[1040] = 25'b0011100001001000010111001;
      square_table[1041] = 25'b0011100000111111000010011;
      square_table[1042] = 25'b0011100000110101101110000;
      square_table[1043] = 25'b0011100000101100011010011;
      square_table[1044] = 25'b0011100000100011000111010;
      square_table[1045] = 25'b0011100000011001110100110;
      square_table[1046] = 25'b0011100000010000100010110;
      square_table[1047] = 25'b0011100000000111010001010;
      square_table[1048] = 25'b0011011111111110000000101;
      square_table[1049] = 25'b0011011111110100110000010;
      square_table[1050] = 25'b0011011111101011100000101;
      square_table[1051] = 25'b0011011111100010010001101;
      square_table[1052] = 25'b0011011111011001000011000;
      square_table[1053] = 25'b0011011111001111110101001;
      square_table[1054] = 25'b0011011111000110100111101;
      square_table[1055] = 25'b0011011110111101011010111;
      square_table[1056] = 25'b0011011110110100001110110;
      square_table[1057] = 25'b0011011110101011000011000;
      square_table[1058] = 25'b0011011110100001110111111;
      square_table[1059] = 25'b0011011110011000101101011;
      square_table[1060] = 25'b0011011110001111100011011;
      square_table[1061] = 25'b0011011110000110011010000;
      square_table[1062] = 25'b0011011101111101010001000;
      square_table[1063] = 25'b0011011101110100001000110;
      square_table[1064] = 25'b0011011101101011000001000;
      square_table[1065] = 25'b0011011101100001111010000;
      square_table[1066] = 25'b0011011101011000110011010;
      square_table[1067] = 25'b0011011101001111101101010;
      square_table[1068] = 25'b0011011101000110101000000;
      square_table[1069] = 25'b0011011100111101100011000;
      square_table[1070] = 25'b0011011100110100011110101;
      square_table[1071] = 25'b0011011100101011011010111;
      square_table[1072] = 25'b0011011100100010010111101;
      square_table[1073] = 25'b0011011100011001010101000;
      square_table[1074] = 25'b0011011100010000010010110;
      square_table[1075] = 25'b0011011100000111010001001;
      square_table[1076] = 25'b0011011011111110010000010;
      square_table[1077] = 25'b0011011011110101001111101;
      square_table[1078] = 25'b0011011011101100001111110;
      square_table[1079] = 25'b0011011011100011010000011;
      square_table[1080] = 25'b0011011011011010010001110;
      square_table[1081] = 25'b0011011011010001010011011;
      square_table[1082] = 25'b0011011011001000010101110;
      square_table[1083] = 25'b0011011010111111011000101;
      square_table[1084] = 25'b0011011010110110011011111;
      square_table[1085] = 25'b0011011010101101100000000;
      square_table[1086] = 25'b0011011010100100100100011;
      square_table[1087] = 25'b0011011010011011101001011;
      square_table[1088] = 25'b0011011010010010101111001;
      square_table[1089] = 25'b0011011010001001110101001;
      square_table[1090] = 25'b0011011010000000111011111;
      square_table[1091] = 25'b0011011001111000000011001;
      square_table[1092] = 25'b0011011001101111001010111;
      square_table[1093] = 25'b0011011001100110010011001;
      square_table[1094] = 25'b0011011001011101011100000;
      square_table[1095] = 25'b0011011001010100100101010;
      square_table[1096] = 25'b0011011001001011101111010;
      square_table[1097] = 25'b0011011001000010111001101;
      square_table[1098] = 25'b0011011000111010000100110;
      square_table[1099] = 25'b0011011000110001010000010;
      square_table[1100] = 25'b0011011000101000011100011;
      square_table[1101] = 25'b0011011000011111101001000;
      square_table[1102] = 25'b0011011000010110110110001;
      square_table[1103] = 25'b0011011000001110000011111;
      square_table[1104] = 25'b0011011000000101010010000;
      square_table[1105] = 25'b0011010111111100100000110;
      square_table[1106] = 25'b0011010111110011110000001;
      square_table[1107] = 25'b0011010111101010111111111;
      square_table[1108] = 25'b0011010111100010010000011;
      square_table[1109] = 25'b0011010111011001100001001;
      square_table[1110] = 25'b0011010111010000110010101;
      square_table[1111] = 25'b0011010111001000000100101;
      square_table[1112] = 25'b0011010110111111010111001;
      square_table[1113] = 25'b0011010110110110101010000;
      square_table[1114] = 25'b0011010110101101111101100;
      square_table[1115] = 25'b0011010110100101010001101;
      square_table[1116] = 25'b0011010110011100100110010;
      square_table[1117] = 25'b0011010110010011111011011;
      square_table[1118] = 25'b0011010110001011010001000;
      square_table[1119] = 25'b0011010110000010100111001;
      square_table[1120] = 25'b0011010101111001111101110;
      square_table[1121] = 25'b0011010101110001010101001;
      square_table[1122] = 25'b0011010101101000101100111;
      square_table[1123] = 25'b0011010101100000000101001;
      square_table[1124] = 25'b0011010101010111011101111;
      square_table[1125] = 25'b0011010101001110110111010;
      square_table[1126] = 25'b0011010101000110010001000;
      square_table[1127] = 25'b0011010100111101101011011;
      square_table[1128] = 25'b0011010100110101000110011;
      square_table[1129] = 25'b0011010100101100100001101;
      square_table[1130] = 25'b0011010100100011111101100;
      square_table[1131] = 25'b0011010100011011011001111;
      square_table[1132] = 25'b0011010100010010110111000;
      square_table[1133] = 25'b0011010100001010010100011;
      square_table[1134] = 25'b0011010100000001110010010;
      square_table[1135] = 25'b0011010011111001010000110;
      square_table[1136] = 25'b0011010011110000101111111;
      square_table[1137] = 25'b0011010011101000001111011;
      square_table[1138] = 25'b0011010011011111101111011;
      square_table[1139] = 25'b0011010011010111001111111;
      square_table[1140] = 25'b0011010011001110110000111;
      square_table[1141] = 25'b0011010011000110010010011;
      square_table[1142] = 25'b0011010010111101110100100;
      square_table[1143] = 25'b0011010010110101010111000;
      square_table[1144] = 25'b0011010010101100111010001;
      square_table[1145] = 25'b0011010010100100011101110;
      square_table[1146] = 25'b0011010010011100000001111;
      square_table[1147] = 25'b0011010010010011100110100;
      square_table[1148] = 25'b0011010010001011001011100;
      square_table[1149] = 25'b0011010010000010110001001;
      square_table[1150] = 25'b0011010001111010010111011;
      square_table[1151] = 25'b0011010001110001111101111;
      square_table[1152] = 25'b0011010001101001100101001;
      square_table[1153] = 25'b0011010001100001001100101;
      square_table[1154] = 25'b0011010001011000110100110;
      square_table[1155] = 25'b0011010001010000011101100;
      square_table[1156] = 25'b0011010001001000000110101;
      square_table[1157] = 25'b0011010000111111110000010;
      square_table[1158] = 25'b0011010000110111011010011;
      square_table[1159] = 25'b0011010000101111000101000;
      square_table[1160] = 25'b0011010000100110110000010;
      square_table[1161] = 25'b0011010000011110011011110;
      square_table[1162] = 25'b0011010000010110000111111;
      square_table[1163] = 25'b0011010000001101110100101;
      square_table[1164] = 25'b0011010000000101100001101;
      square_table[1165] = 25'b0011001111111101001111010;
      square_table[1166] = 25'b0011001111110100111101011;
      square_table[1167] = 25'b0011001111101100101100001;
      square_table[1168] = 25'b0011001111100100011011000;
      square_table[1169] = 25'b0011001111011100001010101;
      square_table[1170] = 25'b0011001111010011111010110;
      square_table[1171] = 25'b0011001111001011101011010;
      square_table[1172] = 25'b0011001111000011011100100;
      square_table[1173] = 25'b0011001110111011001110000;
      square_table[1174] = 25'b0011001110110011000000001;
      square_table[1175] = 25'b0011001110101010110010101;
      square_table[1176] = 25'b0011001110100010100101110;
      square_table[1177] = 25'b0011001110011010011001001;
      square_table[1178] = 25'b0011001110010010001101001;
      square_table[1179] = 25'b0011001110001010000001101;
      square_table[1180] = 25'b0011001110000001110110101;
      square_table[1181] = 25'b0011001101111001101100001;
      square_table[1182] = 25'b0011001101110001100010000;
      square_table[1183] = 25'b0011001101101001011000100;
      square_table[1184] = 25'b0011001101100001001111011;
      square_table[1185] = 25'b0011001101011001000110110;
      square_table[1186] = 25'b0011001101010000111110101;
      square_table[1187] = 25'b0011001101001000110111000;
      square_table[1188] = 25'b0011001101000000101111111;
      square_table[1189] = 25'b0011001100111000101001010;
      square_table[1190] = 25'b0011001100110000100011000;
      square_table[1191] = 25'b0011001100101000011101010;
      square_table[1192] = 25'b0011001100100000011000000;
      square_table[1193] = 25'b0011001100011000010011010;
      square_table[1194] = 25'b0011001100010000001111000;
      square_table[1195] = 25'b0011001100001000001011010;
      square_table[1196] = 25'b0011001100000000001000000;
      square_table[1197] = 25'b0011001011111000000101001;
      square_table[1198] = 25'b0011001011110000000010110;
      square_table[1199] = 25'b0011001011101000000000111;
      square_table[1200] = 25'b0011001011011111111111011;
      square_table[1201] = 25'b0011001011010111111110100;
      square_table[1202] = 25'b0011001011001111111110000;
      square_table[1203] = 25'b0011001011000111111110000;
      square_table[1204] = 25'b0011001010111111111110100;
      square_table[1205] = 25'b0011001010110111111111011;
      square_table[1206] = 25'b0011001010110000000000111;
      square_table[1207] = 25'b0011001010101000000010110;
      square_table[1208] = 25'b0011001010100000000101001;
      square_table[1209] = 25'b0011001010011000000111111;
      square_table[1210] = 25'b0011001010010000001011010;
      square_table[1211] = 25'b0011001010001000001111000;
      square_table[1212] = 25'b0011001010000000010011010;
      square_table[1213] = 25'b0011001001111000010111111;
      square_table[1214] = 25'b0011001001110000011101001;
      square_table[1215] = 25'b0011001001101000100010101;
      square_table[1216] = 25'b0011001001100000101000110;
      square_table[1217] = 25'b0011001001011000101111010;
      square_table[1218] = 25'b0011001001010000110110011;
      square_table[1219] = 25'b0011001001001000111101111;
      square_table[1220] = 25'b0011001001000001000101110;
      square_table[1221] = 25'b0011001000111001001110001;
      square_table[1222] = 25'b0011001000110001010111001;
      square_table[1223] = 25'b0011001000101001100000011;
      square_table[1224] = 25'b0011001000100001101010010;
      square_table[1225] = 25'b0011001000011001110100100;
      square_table[1226] = 25'b0011001000010001111111001;
      square_table[1227] = 25'b0011001000001010001010011;
      square_table[1228] = 25'b0011001000000010010110000;
      square_table[1229] = 25'b0011000111111010100010000;
      square_table[1230] = 25'b0011000111110010101110101;
      square_table[1231] = 25'b0011000111101010111011101;
      square_table[1232] = 25'b0011000111100011001001000;
      square_table[1233] = 25'b0011000111011011010111001;
      square_table[1234] = 25'b0011000111010011100101100;
      square_table[1235] = 25'b0011000111001011110100010;
      square_table[1236] = 25'b0011000111000100000011100;
      square_table[1237] = 25'b0011000110111100010011010;
      square_table[1238] = 25'b0011000110110100100011100;
      square_table[1239] = 25'b0011000110101100110100000;
      square_table[1240] = 25'b0011000110100101000101001;
      square_table[1241] = 25'b0011000110011101010110110;
      square_table[1242] = 25'b0011000110010101101000110;
      square_table[1243] = 25'b0011000110001101111011001;
      square_table[1244] = 25'b0011000110000110001110001;
      square_table[1245] = 25'b0011000101111110100001011;
      square_table[1246] = 25'b0011000101110110110101001;
      square_table[1247] = 25'b0011000101101111001001100;
      square_table[1248] = 25'b0011000101100111011110001;
      square_table[1249] = 25'b0011000101011111110011010;
      square_table[1250] = 25'b0011000101011000001000111;
      square_table[1251] = 25'b0011000101010000011110111;
      square_table[1252] = 25'b0011000101001000110101011;
      square_table[1253] = 25'b0011000101000001001100001;
      square_table[1254] = 25'b0011000100111001100011101;
      square_table[1255] = 25'b0011000100110001111011100;
      square_table[1256] = 25'b0011000100101010010011101;
      square_table[1257] = 25'b0011000100100010101100010;
      square_table[1258] = 25'b0011000100011011000101100;
      square_table[1259] = 25'b0011000100010011011111000;
      square_table[1260] = 25'b0011000100001011111001000;
      square_table[1261] = 25'b0011000100000100010011100;
      square_table[1262] = 25'b0011000011111100101110011;
      square_table[1263] = 25'b0011000011110101001001110;
      square_table[1264] = 25'b0011000011101101100101100;
      square_table[1265] = 25'b0011000011100110000001110;
      square_table[1266] = 25'b0011000011011110011110011;
      square_table[1267] = 25'b0011000011010110111011100;
      square_table[1268] = 25'b0011000011001111011001000;
      square_table[1269] = 25'b0011000011000111110111000;
      square_table[1270] = 25'b0011000011000000010101011;
      square_table[1271] = 25'b0011000010111000110100010;
      square_table[1272] = 25'b0011000010110001010011011;
      square_table[1273] = 25'b0011000010101001110011001;
      square_table[1274] = 25'b0011000010100010010011001;
      square_table[1275] = 25'b0011000010011010110011111;
      square_table[1276] = 25'b0011000010010011010100110;
      square_table[1277] = 25'b0011000010001011110110010;
      square_table[1278] = 25'b0011000010000100011000001;
      square_table[1279] = 25'b0011000001111100111010011;
      square_table[1280] = 25'b0011000001110101011101001;
      square_table[1281] = 25'b0011000001101110000000010;
      square_table[1282] = 25'b0011000001100110100011111;
      square_table[1283] = 25'b0011000001011111000111111;
      square_table[1284] = 25'b0011000001010111101100010;
      square_table[1285] = 25'b0011000001010000010001001;
      square_table[1286] = 25'b0011000001001000110110100;
      square_table[1287] = 25'b0011000001000001011100010;
      square_table[1288] = 25'b0011000000111010000010010;
      square_table[1289] = 25'b0011000000110010101001000;
      square_table[1290] = 25'b0011000000101011001111111;
      square_table[1291] = 25'b0011000000100011110111011;
      square_table[1292] = 25'b0011000000011100011111010;
      square_table[1293] = 25'b0011000000010101000111100;
      square_table[1294] = 25'b0011000000001101110000001;
      square_table[1295] = 25'b0011000000000110011001010;
      square_table[1296] = 25'b0010111111111111000010110;
      square_table[1297] = 25'b0010111111110111101100110;
      square_table[1298] = 25'b0010111111110000010111001;
      square_table[1299] = 25'b0010111111101001000010000;
      square_table[1300] = 25'b0010111111100001101101010;
      square_table[1301] = 25'b0010111111011010011000110;
      square_table[1302] = 25'b0010111111010011000101000;
      square_table[1303] = 25'b0010111111001011110001011;
      square_table[1304] = 25'b0010111111000100011110011;
      square_table[1305] = 25'b0010111110111101001011110;
      square_table[1306] = 25'b0010111110110101111001011;
      square_table[1307] = 25'b0010111110101110100111101;
      square_table[1308] = 25'b0010111110100111010110001;
      square_table[1309] = 25'b0010111110100000000101001;
      square_table[1310] = 25'b0010111110011000110100100;
      square_table[1311] = 25'b0010111110010001100100011;
      square_table[1312] = 25'b0010111110001010010100100;
      square_table[1313] = 25'b0010111110000011000101001;
      square_table[1314] = 25'b0010111101111011110110010;
      square_table[1315] = 25'b0010111101110100100111101;
      square_table[1316] = 25'b0010111101101101011001100;
      square_table[1317] = 25'b0010111101100110001011111;
      square_table[1318] = 25'b0010111101011110111110100;
      square_table[1319] = 25'b0010111101010111110001101;
      square_table[1320] = 25'b0010111101010000100101010;
      square_table[1321] = 25'b0010111101001001011001001;
      square_table[1322] = 25'b0010111101000010001101101;
      square_table[1323] = 25'b0010111100111011000010010;
      square_table[1324] = 25'b0010111100110011110111011;
      square_table[1325] = 25'b0010111100101100101101000;
      square_table[1326] = 25'b0010111100100101100011000;
      square_table[1327] = 25'b0010111100011110011001011;
      square_table[1328] = 25'b0010111100010111010000001;
      square_table[1329] = 25'b0010111100010000000111011;
      square_table[1330] = 25'b0010111100001000111110111;
      square_table[1331] = 25'b0010111100000001110111000;
      square_table[1332] = 25'b0010111011111010101111100;
      square_table[1333] = 25'b0010111011110011101000010;
      square_table[1334] = 25'b0010111011101100100001100;
      square_table[1335] = 25'b0010111011100101011011000;
      square_table[1336] = 25'b0010111011011110010101001;
      square_table[1337] = 25'b0010111011010111001111100;
      square_table[1338] = 25'b0010111011010000001010010;
      square_table[1339] = 25'b0010111011001001000101100;
      square_table[1340] = 25'b0010111011000010000001010;
      square_table[1341] = 25'b0010111010111010111101010;
      square_table[1342] = 25'b0010111010110011111001101;
      square_table[1343] = 25'b0010111010101100110110100;
      square_table[1344] = 25'b0010111010100101110011110;
      square_table[1345] = 25'b0010111010011110110001011;
      square_table[1346] = 25'b0010111010010111101111100;
      square_table[1347] = 25'b0010111010010000101101110;
      square_table[1348] = 25'b0010111010001001101100101;
      square_table[1349] = 25'b0010111010000010101100000;
      square_table[1350] = 25'b0010111001111011101011100;
      square_table[1351] = 25'b0010111001110100101011100;
      square_table[1352] = 25'b0010111001101101101011111;
      square_table[1353] = 25'b0010111001100110101100110;
      square_table[1354] = 25'b0010111001011111101101111;
      square_table[1355] = 25'b0010111001011000101111100;
      square_table[1356] = 25'b0010111001010001110001100;
      square_table[1357] = 25'b0010111001001010110011111;
      square_table[1358] = 25'b0010111001000011110110101;
      square_table[1359] = 25'b0010111000111100111001110;
      square_table[1360] = 25'b0010111000110101111101011;
      square_table[1361] = 25'b0010111000101111000001010;
      square_table[1362] = 25'b0010111000101000000101101;
      square_table[1363] = 25'b0010111000100001001010011;
      square_table[1364] = 25'b0010111000011010001111100;
      square_table[1365] = 25'b0010111000010011010101000;
      square_table[1366] = 25'b0010111000001100011010111;
      square_table[1367] = 25'b0010111000000101100001001;
      square_table[1368] = 25'b0010110111111110100111110;
      square_table[1369] = 25'b0010110111110111101110111;
      square_table[1370] = 25'b0010110111110000110110011;
      square_table[1371] = 25'b0010110111101001111110001;
      square_table[1372] = 25'b0010110111100011000110011;
      square_table[1373] = 25'b0010110111011100001111000;
      square_table[1374] = 25'b0010110111010101010111111;
      square_table[1375] = 25'b0010110111001110100001010;
      square_table[1376] = 25'b0010110111000111101011000;
      square_table[1377] = 25'b0010110111000000110101001;
      square_table[1378] = 25'b0010110110111001111111110;
      square_table[1379] = 25'b0010110110110011001010101;
      square_table[1380] = 25'b0010110110101100010101111;
      square_table[1381] = 25'b0010110110100101100001101;
      square_table[1382] = 25'b0010110110011110101101100;
      square_table[1383] = 25'b0010110110010111111010001;
      square_table[1384] = 25'b0010110110010001000110110;
      square_table[1385] = 25'b0010110110001010010100000;
      square_table[1386] = 25'b0010110110000011100001101;
      square_table[1387] = 25'b0010110101111100101111100;
      square_table[1388] = 25'b0010110101110101111101111;
      square_table[1389] = 25'b0010110101101111001100101;
      square_table[1390] = 25'b0010110101101000011011101;
      square_table[1391] = 25'b0010110101100001101011001;
      square_table[1392] = 25'b0010110101011010111010111;
      square_table[1393] = 25'b0010110101010100001011010;
      square_table[1394] = 25'b0010110101001101011011110;
      square_table[1395] = 25'b0010110101000110101100110;
      square_table[1396] = 25'b0010110100111111111110001;
      square_table[1397] = 25'b0010110100111001001111111;
      square_table[1398] = 25'b0010110100110010100001111;
      square_table[1399] = 25'b0010110100101011110100100;
      square_table[1400] = 25'b0010110100100101000111001;
      square_table[1401] = 25'b0010110100011110011010100;
      square_table[1402] = 25'b0010110100010111101110000;
      square_table[1403] = 25'b0010110100010001000010000;
      square_table[1404] = 25'b0010110100001010010110011;
      square_table[1405] = 25'b0010110100000011101011000;
      square_table[1406] = 25'b0010110011111101000000001;
      square_table[1407] = 25'b0010110011110110010101101;
      square_table[1408] = 25'b0010110011101111101011011;
      square_table[1409] = 25'b0010110011101001000001101;
      square_table[1410] = 25'b0010110011100010011000001;
      square_table[1411] = 25'b0010110011011011101111000;
      square_table[1412] = 25'b0010110011010101000110010;
      square_table[1413] = 25'b0010110011001110011110000;
      square_table[1414] = 25'b0010110011000111110110000;
      square_table[1415] = 25'b0010110011000001001110011;
      square_table[1416] = 25'b0010110010111010100111010;
      square_table[1417] = 25'b0010110010110100000000011;
      square_table[1418] = 25'b0010110010101101011001111;
      square_table[1419] = 25'b0010110010100110110011101;
      square_table[1420] = 25'b0010110010100000001101111;
      square_table[1421] = 25'b0010110010011001101000100;
      square_table[1422] = 25'b0010110010010011000011011;
      square_table[1423] = 25'b0010110010001100011110101;
      square_table[1424] = 25'b0010110010000101111010011;
      square_table[1425] = 25'b0010110001111111010110011;
      square_table[1426] = 25'b0010110001111000110010110;
      square_table[1427] = 25'b0010110001110010001111101;
      square_table[1428] = 25'b0010110001101011101100110;
      square_table[1429] = 25'b0010110001100101001010010;
      square_table[1430] = 25'b0010110001011110101000001;
      square_table[1431] = 25'b0010110001011000000110010;
      square_table[1432] = 25'b0010110001010001100100111;
      square_table[1433] = 25'b0010110001001011000011110;
      square_table[1434] = 25'b0010110001000100100011000;
      square_table[1435] = 25'b0010110000111110000010110;
      square_table[1436] = 25'b0010110000110111100010110;
      square_table[1437] = 25'b0010110000110001000011001;
      square_table[1438] = 25'b0010110000101010100011111;
      square_table[1439] = 25'b0010110000100100000101000;
      square_table[1440] = 25'b0010110000011101100110011;
      square_table[1441] = 25'b0010110000010111001000001;
      square_table[1442] = 25'b0010110000010000101010010;
      square_table[1443] = 25'b0010110000001010001100111;
      square_table[1444] = 25'b0010110000000011101111101;
      square_table[1445] = 25'b0010101111111101010010111;
      square_table[1446] = 25'b0010101111110110110110011;
      square_table[1447] = 25'b0010101111110000011010010;
      square_table[1448] = 25'b0010101111101001111110101;
      square_table[1449] = 25'b0010101111100011100011010;
      square_table[1450] = 25'b0010101111011101001000010;
      square_table[1451] = 25'b0010101111010110101101101;
      square_table[1452] = 25'b0010101111010000010011010;
      square_table[1453] = 25'b0010101111001001111001011;
      square_table[1454] = 25'b0010101111000011011111110;
      square_table[1455] = 25'b0010101110111101000110100;
      square_table[1456] = 25'b0010101110110110101101100;
      square_table[1457] = 25'b0010101110110000010100111;
      square_table[1458] = 25'b0010101110101001111100110;
      square_table[1459] = 25'b0010101110100011100101000;
      square_table[1460] = 25'b0010101110011101001101011;
      square_table[1461] = 25'b0010101110010110110110010;
      square_table[1462] = 25'b0010101110010000011111011;
      square_table[1463] = 25'b0010101110001010001001000;
      square_table[1464] = 25'b0010101110000011110010111;
      square_table[1465] = 25'b0010101101111101011101001;
      square_table[1466] = 25'b0010101101110111000111101;
      square_table[1467] = 25'b0010101101110000110010100;
      square_table[1468] = 25'b0010101101101010011101111;
      square_table[1469] = 25'b0010101101100100001001011;
      square_table[1470] = 25'b0010101101011101110101011;
      square_table[1471] = 25'b0010101101010111100001101;
      square_table[1472] = 25'b0010101101010001001110010;
      square_table[1473] = 25'b0010101101001010111011010;
      square_table[1474] = 25'b0010101101000100101000100;
      square_table[1475] = 25'b0010101100111110010110010;
      square_table[1476] = 25'b0010101100111000000100010;
      square_table[1477] = 25'b0010101100110001110010101;
      square_table[1478] = 25'b0010101100101011100001010;
      square_table[1479] = 25'b0010101100100101010000011;
      square_table[1480] = 25'b0010101100011110111111110;
      square_table[1481] = 25'b0010101100011000101111100;
      square_table[1482] = 25'b0010101100010010011111100;
      square_table[1483] = 25'b0010101100001100010000000;
      square_table[1484] = 25'b0010101100000110000000101;
      square_table[1485] = 25'b0010101011111111110001110;
      square_table[1486] = 25'b0010101011111001100011001;
      square_table[1487] = 25'b0010101011110011010100111;
      square_table[1488] = 25'b0010101011101101000111000;
      square_table[1489] = 25'b0010101011100110111001011;
      square_table[1490] = 25'b0010101011100000101100001;
      square_table[1491] = 25'b0010101011011010011111010;
      square_table[1492] = 25'b0010101011010100010010110;
      square_table[1493] = 25'b0010101011001110000110100;
      square_table[1494] = 25'b0010101011000111111010101;
      square_table[1495] = 25'b0010101011000001101111001;
      square_table[1496] = 25'b0010101010111011100011111;
      square_table[1497] = 25'b0010101010110101011001000;
      square_table[1498] = 25'b0010101010101111001110011;
      square_table[1499] = 25'b0010101010101001000100001;
      square_table[1500] = 25'b0010101010100010111010011;
      square_table[1501] = 25'b0010101010011100110000110;
      square_table[1502] = 25'b0010101010010110100111101;
      square_table[1503] = 25'b0010101010010000011110110;
      square_table[1504] = 25'b0010101010001010010110000;
      square_table[1505] = 25'b0010101010000100001101110;
      square_table[1506] = 25'b0010101001111110000110000;
      square_table[1507] = 25'b0010101001110111111110011;
      square_table[1508] = 25'b0010101001110001110111001;
      square_table[1509] = 25'b0010101001101011110000010;
      square_table[1510] = 25'b0010101001100101101001101;
      square_table[1511] = 25'b0010101001011111100011100;
      square_table[1512] = 25'b0010101001011001011101101;
      square_table[1513] = 25'b0010101001010011011000000;
      square_table[1514] = 25'b0010101001001101010010110;
      square_table[1515] = 25'b0010101001000111001101110;
      square_table[1516] = 25'b0010101001000001001001001;
      square_table[1517] = 25'b0010101000111011000100111;
      square_table[1518] = 25'b0010101000110101000001000;
      square_table[1519] = 25'b0010101000101110111101010;
      square_table[1520] = 25'b0010101000101000111010000;
      square_table[1521] = 25'b0010101000100010110111001;
      square_table[1522] = 25'b0010101000011100110100011;
      square_table[1523] = 25'b0010101000010110110010000;
      square_table[1524] = 25'b0010101000010000110000000;
      square_table[1525] = 25'b0010101000001010101110011;
      square_table[1526] = 25'b0010101000000100101101000;
      square_table[1527] = 25'b0010100111111110101100001;
      square_table[1528] = 25'b0010100111111000101011011;
      square_table[1529] = 25'b0010100111110010101010111;
      square_table[1530] = 25'b0010100111101100101010111;
      square_table[1531] = 25'b0010100111100110101011001;
      square_table[1532] = 25'b0010100111100000101011110;
      square_table[1533] = 25'b0010100111011010101100110;
      square_table[1534] = 25'b0010100111010100101101111;
      square_table[1535] = 25'b0010100111001110101111011;
      square_table[1536] = 25'b0010100111001000110001010;
      square_table[1537] = 25'b0010100111000010110011100;
      square_table[1538] = 25'b0010100110111100110110000;
      square_table[1539] = 25'b0010100110110110111000110;
      square_table[1540] = 25'b0010100110110000111011111;
      square_table[1541] = 25'b0010100110101010111111011;
      square_table[1542] = 25'b0010100110100101000011001;
      square_table[1543] = 25'b0010100110011111000111010;
      square_table[1544] = 25'b0010100110011001001011101;
      square_table[1545] = 25'b0010100110010011010000011;
      square_table[1546] = 25'b0010100110001101010101100;
      square_table[1547] = 25'b0010100110000111011010110;
      square_table[1548] = 25'b0010100110000001100000100;
      square_table[1549] = 25'b0010100101111011100110011;
      square_table[1550] = 25'b0010100101110101101100110;
      square_table[1551] = 25'b0010100101101111110011100;
      square_table[1552] = 25'b0010100101101001111010010;
      square_table[1553] = 25'b0010100101100100000001101;
      square_table[1554] = 25'b0010100101011110001001001;
      square_table[1555] = 25'b0010100101011000010001001;
      square_table[1556] = 25'b0010100101010010011001010;
      square_table[1557] = 25'b0010100101001100100001110;
      square_table[1558] = 25'b0010100101000110101010101;
      square_table[1559] = 25'b0010100101000000110011110;
      square_table[1560] = 25'b0010100100111010111101010;
      square_table[1561] = 25'b0010100100110101000111000;
      square_table[1562] = 25'b0010100100101111010001000;
      square_table[1563] = 25'b0010100100101001011011011;
      square_table[1564] = 25'b0010100100100011100110000;
      square_table[1565] = 25'b0010100100011101110001000;
      square_table[1566] = 25'b0010100100010111111100010;
      square_table[1567] = 25'b0010100100010010000111111;
      square_table[1568] = 25'b0010100100001100010011110;
      square_table[1569] = 25'b0010100100000110100000001;
      square_table[1570] = 25'b0010100100000000101100101;
      square_table[1571] = 25'b0010100011111010111001100;
      square_table[1572] = 25'b0010100011110101000110101;
      square_table[1573] = 25'b0010100011101111010100001;
      square_table[1574] = 25'b0010100011101001100001111;
      square_table[1575] = 25'b0010100011100011101111111;
      square_table[1576] = 25'b0010100011011101111110010;
      square_table[1577] = 25'b0010100011011000001101000;
      square_table[1578] = 25'b0010100011010010011100000;
      square_table[1579] = 25'b0010100011001100101011010;
      square_table[1580] = 25'b0010100011000110111010111;
      square_table[1581] = 25'b0010100011000001001010111;
      square_table[1582] = 25'b0010100010111011011011000;
      square_table[1583] = 25'b0010100010110101101011100;
      square_table[1584] = 25'b0010100010101111111100010;
      square_table[1585] = 25'b0010100010101010001101100;
      square_table[1586] = 25'b0010100010100100011110111;
      square_table[1587] = 25'b0010100010011110110000101;
      square_table[1588] = 25'b0010100010011001000010101;
      square_table[1589] = 25'b0010100010010011010100111;
      square_table[1590] = 25'b0010100010001101100111101;
      square_table[1591] = 25'b0010100010000111111010100;
      square_table[1592] = 25'b0010100010000010001101110;
      square_table[1593] = 25'b0010100001111100100001010;
      square_table[1594] = 25'b0010100001110110110101001;
      square_table[1595] = 25'b0010100001110001001001010;
      square_table[1596] = 25'b0010100001101011011101101;
      square_table[1597] = 25'b0010100001100101110010011;
      square_table[1598] = 25'b0010100001100000000111011;
      square_table[1599] = 25'b0010100001011010011100110;
      square_table[1600] = 25'b0010100001010100110010011;
      square_table[1601] = 25'b0010100001001111001000011;
      square_table[1602] = 25'b0010100001001001011110101;
      square_table[1603] = 25'b0010100001000011110101001;
      square_table[1604] = 25'b0010100000111110001011111;
      square_table[1605] = 25'b0010100000111000100011000;
      square_table[1606] = 25'b0010100000110010111010011;
      square_table[1607] = 25'b0010100000101101010010000;
      square_table[1608] = 25'b0010100000100111101010001;
      square_table[1609] = 25'b0010100000100010000010100;
      square_table[1610] = 25'b0010100000011100011011000;
      square_table[1611] = 25'b0010100000010110110011111;
      square_table[1612] = 25'b0010100000010001001101000;
      square_table[1613] = 25'b0010100000001011100110101;
      square_table[1614] = 25'b0010100000000110000000011;
      square_table[1615] = 25'b0010100000000000011010011;
      square_table[1616] = 25'b0010011111111010110100101;
      square_table[1617] = 25'b0010011111110101001111011;
      square_table[1618] = 25'b0010011111101111101010011;
      square_table[1619] = 25'b0010011111101010000101100;
      square_table[1620] = 25'b0010011111100100100001001;
      square_table[1621] = 25'b0010011111011110111100111;
      square_table[1622] = 25'b0010011111011001011001000;
      square_table[1623] = 25'b0010011111010011110101100;
      square_table[1624] = 25'b0010011111001110010010000;
      square_table[1625] = 25'b0010011111001000101111000;
      square_table[1626] = 25'b0010011111000011001100011;
      square_table[1627] = 25'b0010011110111101101001111;
      square_table[1628] = 25'b0010011110111000000111110;
      square_table[1629] = 25'b0010011110110010100101111;
      square_table[1630] = 25'b0010011110101101000100010;
      square_table[1631] = 25'b0010011110100111100011000;
      square_table[1632] = 25'b0010011110100010000010000;
      square_table[1633] = 25'b0010011110011100100001010;
      square_table[1634] = 25'b0010011110010111000000111;
      square_table[1635] = 25'b0010011110010001100000110;
      square_table[1636] = 25'b0010011110001100000000111;
      square_table[1637] = 25'b0010011110000110100001011;
      square_table[1638] = 25'b0010011110000001000010000;
      square_table[1639] = 25'b0010011101111011100011000;
      square_table[1640] = 25'b0010011101110110000100010;
      square_table[1641] = 25'b0010011101110000100101111;
      square_table[1642] = 25'b0010011101101011000111110;
      square_table[1643] = 25'b0010011101100101101001111;
      square_table[1644] = 25'b0010011101100000001100011;
      square_table[1645] = 25'b0010011101011010101111000;
      square_table[1646] = 25'b0010011101010101010010000;
      square_table[1647] = 25'b0010011101001111110101011;
      square_table[1648] = 25'b0010011101001010011000111;
      square_table[1649] = 25'b0010011101000100111100110;
      square_table[1650] = 25'b0010011100111111100000111;
      square_table[1651] = 25'b0010011100111010000101010;
      square_table[1652] = 25'b0010011100110100101001111;
      square_table[1653] = 25'b0010011100101111001111000;
      square_table[1654] = 25'b0010011100101001110100001;
      square_table[1655] = 25'b0010011100100100011001110;
      square_table[1656] = 25'b0010011100011110111111100;
      square_table[1657] = 25'b0010011100011001100101101;
      square_table[1658] = 25'b0010011100010100001011111;
      square_table[1659] = 25'b0010011100001110110010101;
      square_table[1660] = 25'b0010011100001001011001101;
      square_table[1661] = 25'b0010011100000100000000110;
      square_table[1662] = 25'b0010011011111110101000010;
      square_table[1663] = 25'b0010011011111001010000000;
      square_table[1664] = 25'b0010011011110011111000000;
      square_table[1665] = 25'b0010011011101110100000011;
      square_table[1666] = 25'b0010011011101001001001000;
      square_table[1667] = 25'b0010011011100011110010000;
      square_table[1668] = 25'b0010011011011110011011000;
      square_table[1669] = 25'b0010011011011001000100100;
      square_table[1670] = 25'b0010011011010011101110010;
      square_table[1671] = 25'b0010011011001110011000001;
      square_table[1672] = 25'b0010011011001001000010100;
      square_table[1673] = 25'b0010011011000011101101000;
      square_table[1674] = 25'b0010011010111110010111111;
      square_table[1675] = 25'b0010011010111001000011000;
      square_table[1676] = 25'b0010011010110011101110010;
      square_table[1677] = 25'b0010011010101110011001111;
      square_table[1678] = 25'b0010011010101001000101111;
      square_table[1679] = 25'b0010011010100011110010000;
      square_table[1680] = 25'b0010011010011110011110100;
      square_table[1681] = 25'b0010011010011001001011010;
      square_table[1682] = 25'b0010011010010011111000001;
      square_table[1683] = 25'b0010011010001110100101100;
      square_table[1684] = 25'b0010011010001001010011000;
      square_table[1685] = 25'b0010011010000100000000110;
      square_table[1686] = 25'b0010011001111110101110111;
      square_table[1687] = 25'b0010011001111001011101010;
      square_table[1688] = 25'b0010011001110100001011111;
      square_table[1689] = 25'b0010011001101110111010111;
      square_table[1690] = 25'b0010011001101001101010000;
      square_table[1691] = 25'b0010011001100100011001100;
      square_table[1692] = 25'b0010011001011111001001010;
      square_table[1693] = 25'b0010011001011001111001010;
      square_table[1694] = 25'b0010011001010100101001100;
      square_table[1695] = 25'b0010011001001111011001111;
      square_table[1696] = 25'b0010011001001010001010110;
      square_table[1697] = 25'b0010011001000100111011110;
      square_table[1698] = 25'b0010011000111111101101010;
      square_table[1699] = 25'b0010011000111010011110110;
      square_table[1700] = 25'b0010011000110101010000100;
      square_table[1701] = 25'b0010011000110000000010110;
      square_table[1702] = 25'b0010011000101010110101001;
      square_table[1703] = 25'b0010011000100101100111110;
      square_table[1704] = 25'b0010011000100000011010110;
      square_table[1705] = 25'b0010011000011011001101111;
      square_table[1706] = 25'b0010011000010110000001011;
      square_table[1707] = 25'b0010011000010000110101001;
      square_table[1708] = 25'b0010011000001011101001010;
      square_table[1709] = 25'b0010011000000110011101011;
      square_table[1710] = 25'b0010011000000001010001111;
      square_table[1711] = 25'b0010010111111100000110110;
      square_table[1712] = 25'b0010010111110110111011110;
      square_table[1713] = 25'b0010010111110001110001001;
      square_table[1714] = 25'b0010010111101100100110101;
      square_table[1715] = 25'b0010010111100111011100100;
      square_table[1716] = 25'b0010010111100010010010101;
      square_table[1717] = 25'b0010010111011101001001000;
      square_table[1718] = 25'b0010010111010111111111101;
      square_table[1719] = 25'b0010010111010010110110101;
      square_table[1720] = 25'b0010010111001101101101110;
      square_table[1721] = 25'b0010010111001000100101001;
      square_table[1722] = 25'b0010010111000011011100110;
      square_table[1723] = 25'b0010010110111110010100110;
      square_table[1724] = 25'b0010010110111001001100111;
      square_table[1725] = 25'b0010010110110100000101100;
      square_table[1726] = 25'b0010010110101110111110001;
      square_table[1727] = 25'b0010010110101001110111001;
      square_table[1728] = 25'b0010010110100100110000011;
      square_table[1729] = 25'b0010010110011111101001111;
      square_table[1730] = 25'b0010010110011010100011100;
      square_table[1731] = 25'b0010010110010101011101101;
      square_table[1732] = 25'b0010010110010000011000000;
      square_table[1733] = 25'b0010010110001011010010011;
      square_table[1734] = 25'b0010010110000110001101010;
      square_table[1735] = 25'b0010010110000001001000010;
      square_table[1736] = 25'b0010010101111100000011100;
      square_table[1737] = 25'b0010010101110110111111001;
      square_table[1738] = 25'b0010010101110001111011000;
      square_table[1739] = 25'b0010010101101100110111001;
      square_table[1740] = 25'b0010010101100111110011100;
      square_table[1741] = 25'b0010010101100010110000000;
      square_table[1742] = 25'b0010010101011101101100111;
      square_table[1743] = 25'b0010010101011000101010000;
      square_table[1744] = 25'b0010010101010011100111011;
      square_table[1745] = 25'b0010010101001110100101000;
      square_table[1746] = 25'b0010010101001001100010111;
      square_table[1747] = 25'b0010010101000100100001000;
      square_table[1748] = 25'b0010010100111111011111011;
      square_table[1749] = 25'b0010010100111010011110000;
      square_table[1750] = 25'b0010010100110101011100111;
      square_table[1751] = 25'b0010010100110000011100000;
      square_table[1752] = 25'b0010010100101011011011100;
      square_table[1753] = 25'b0010010100100110011011001;
      square_table[1754] = 25'b0010010100100001011011000;
      square_table[1755] = 25'b0010010100011100011011001;
      square_table[1756] = 25'b0010010100010111011011100;
      square_table[1757] = 25'b0010010100010010011100001;
      square_table[1758] = 25'b0010010100001101011101001;
      square_table[1759] = 25'b0010010100001000011110010;
      square_table[1760] = 25'b0010010100000011011111101;
      square_table[1761] = 25'b0010010011111110100001011;
      square_table[1762] = 25'b0010010011111001100011010;
      square_table[1763] = 25'b0010010011110100100101011;
      square_table[1764] = 25'b0010010011101111100111110;
      square_table[1765] = 25'b0010010011101010101010100;
      square_table[1766] = 25'b0010010011100101101101011;
      square_table[1767] = 25'b0010010011100000110000100;
      square_table[1768] = 25'b0010010011011011110100000;
      square_table[1769] = 25'b0010010011010110110111101;
      square_table[1770] = 25'b0010010011010001111011100;
      square_table[1771] = 25'b0010010011001100111111101;
      square_table[1772] = 25'b0010010011001000000100001;
      square_table[1773] = 25'b0010010011000011001000110;
      square_table[1774] = 25'b0010010010111110001101101;
      square_table[1775] = 25'b0010010010111001010010110;
      square_table[1776] = 25'b0010010010110100011000010;
      square_table[1777] = 25'b0010010010101111011101111;
      square_table[1778] = 25'b0010010010101010100011110;
      square_table[1779] = 25'b0010010010100101101001111;
      square_table[1780] = 25'b0010010010100000110000010;
      square_table[1781] = 25'b0010010010011011110110111;
      square_table[1782] = 25'b0010010010010110111101110;
      square_table[1783] = 25'b0010010010010010000100111;
      square_table[1784] = 25'b0010010010001101001100010;
      square_table[1785] = 25'b0010010010001000010011110;
      square_table[1786] = 25'b0010010010000011011011110;
      square_table[1787] = 25'b0010010001111110100011111;
      square_table[1788] = 25'b0010010001111001101100001;
      square_table[1789] = 25'b0010010001110100110100110;
      square_table[1790] = 25'b0010010001101111111101100;
      square_table[1791] = 25'b0010010001101011000110101;
      square_table[1792] = 25'b0010010001100110010000000;
      square_table[1793] = 25'b0010010001100001011001100;
      square_table[1794] = 25'b0010010001011100100011010;
      square_table[1795] = 25'b0010010001010111101101010;
      square_table[1796] = 25'b0010010001010010110111100;
      square_table[1797] = 25'b0010010001001110000010001;
      square_table[1798] = 25'b0010010001001001001100111;
      square_table[1799] = 25'b0010010001000100010111110;
      square_table[1800] = 25'b0010010000111111100011001;
      square_table[1801] = 25'b0010010000111010101110101;
      square_table[1802] = 25'b0010010000110101111010010;
      square_table[1803] = 25'b0010010000110001000110011;
      square_table[1804] = 25'b0010010000101100010010100;
      square_table[1805] = 25'b0010010000100111011110111;
      square_table[1806] = 25'b0010010000100010101011101;
      square_table[1807] = 25'b0010010000011101111000100;
      square_table[1808] = 25'b0010010000011001000101101;
      square_table[1809] = 25'b0010010000010100010011001;
      square_table[1810] = 25'b0010010000001111100000110;
      square_table[1811] = 25'b0010010000001010101110101;
      square_table[1812] = 25'b0010010000000101111100110;
      square_table[1813] = 25'b0010010000000001001011001;
      square_table[1814] = 25'b0010001111111100011001101;
      square_table[1815] = 25'b0010001111110111101000100;
      square_table[1816] = 25'b0010001111110010110111100;
      square_table[1817] = 25'b0010001111101110000110111;
      square_table[1818] = 25'b0010001111101001010110011;
      square_table[1819] = 25'b0010001111100100100110010;
      square_table[1820] = 25'b0010001111011111110110001;
      square_table[1821] = 25'b0010001111011011000110100;
      square_table[1822] = 25'b0010001111010110010110111;
      square_table[1823] = 25'b0010001111010001100111100;
      square_table[1824] = 25'b0010001111001100111000101;
      square_table[1825] = 25'b0010001111001000001001110;
      square_table[1826] = 25'b0010001111000011011011010;
      square_table[1827] = 25'b0010001110111110101100110;
      square_table[1828] = 25'b0010001110111001111110101;
      square_table[1829] = 25'b0010001110110101010000110;
      square_table[1830] = 25'b0010001110110000100011010;
      square_table[1831] = 25'b0010001110101011110101110;
      square_table[1832] = 25'b0010001110100111001000101;
      square_table[1833] = 25'b0010001110100010011011101;
      square_table[1834] = 25'b0010001110011101101110111;
      square_table[1835] = 25'b0010001110011001000010100;
      square_table[1836] = 25'b0010001110010100010110010;
      square_table[1837] = 25'b0010001110001111101010001;
      square_table[1838] = 25'b0010001110001010111110011;
      square_table[1839] = 25'b0010001110000110010010111;
      square_table[1840] = 25'b0010001110000001100111100;
      square_table[1841] = 25'b0010001101111100111100011;
      square_table[1842] = 25'b0010001101111000010001100;
      square_table[1843] = 25'b0010001101110011100111000;
      square_table[1844] = 25'b0010001101101110111100101;
      square_table[1845] = 25'b0010001101101010010010010;
      square_table[1846] = 25'b0010001101100101101000011;
      square_table[1847] = 25'b0010001101100000111110110;
      square_table[1848] = 25'b0010001101011100010101010;
      square_table[1849] = 25'b0010001101010111101100000;
      square_table[1850] = 25'b0010001101010011000010111;
      square_table[1851] = 25'b0010001101001110011010001;
      square_table[1852] = 25'b0010001101001001110001101;
      square_table[1853] = 25'b0010001101000101001001010;
      square_table[1854] = 25'b0010001101000000100001001;
      square_table[1855] = 25'b0010001100111011111001010;
      square_table[1856] = 25'b0010001100110111010001100;
      square_table[1857] = 25'b0010001100110010101010001;
      square_table[1858] = 25'b0010001100101110000010111;
      square_table[1859] = 25'b0010001100101001011100000;
      square_table[1860] = 25'b0010001100100100110101001;
      square_table[1861] = 25'b0010001100100000001110110;
      square_table[1862] = 25'b0010001100011011101000011;
      square_table[1863] = 25'b0010001100010111000010011;
      square_table[1864] = 25'b0010001100010010011100100;
      square_table[1865] = 25'b0010001100001101110110111;
      square_table[1866] = 25'b0010001100001001010001100;
      square_table[1867] = 25'b0010001100000100101100010;
      square_table[1868] = 25'b0010001100000000000111010;
      square_table[1869] = 25'b0010001011111011100010101;
      square_table[1870] = 25'b0010001011110110111110001;
      square_table[1871] = 25'b0010001011110010011001111;
      square_table[1872] = 25'b0010001011101101110101111;
      square_table[1873] = 25'b0010001011101001010010000;
      square_table[1874] = 25'b0010001011100100101110011;
      square_table[1875] = 25'b0010001011100000001010111;
      square_table[1876] = 25'b0010001011011011100111111;
      square_table[1877] = 25'b0010001011010111000100110;
      square_table[1878] = 25'b0010001011010010100010001;
      square_table[1879] = 25'b0010001011001101111111101;
      square_table[1880] = 25'b0010001011001001011101011;
      square_table[1881] = 25'b0010001011000100111011010;
      square_table[1882] = 25'b0010001011000000011001100;
      square_table[1883] = 25'b0010001010111011110111111;
      square_table[1884] = 25'b0010001010110111010110100;
      square_table[1885] = 25'b0010001010110010110101011;
      square_table[1886] = 25'b0010001010101110010100011;
      square_table[1887] = 25'b0010001010101001110011101;
      square_table[1888] = 25'b0010001010100101010011010;
      square_table[1889] = 25'b0010001010100000110010111;
      square_table[1890] = 25'b0010001010011100010010110;
      square_table[1891] = 25'b0010001010010111110011000;
      square_table[1892] = 25'b0010001010010011010011010;
      square_table[1893] = 25'b0010001010001110110011111;
      square_table[1894] = 25'b0010001010001010010100110;
      square_table[1895] = 25'b0010001010000101110101110;
      square_table[1896] = 25'b0010001010000001010111000;
      square_table[1897] = 25'b0010001001111100111000100;
      square_table[1898] = 25'b0010001001111000011010001;
      square_table[1899] = 25'b0010001001110011111100000;
      square_table[1900] = 25'b0010001001101111011110001;
      square_table[1901] = 25'b0010001001101011000000100;
      square_table[1902] = 25'b0010001001100110100011000;
      square_table[1903] = 25'b0010001001100010000101111;
      square_table[1904] = 25'b0010001001011101101000110;
      square_table[1905] = 25'b0010001001011001001100000;
      square_table[1906] = 25'b0010001001010100101111011;
      square_table[1907] = 25'b0010001001010000010011001;
      square_table[1908] = 25'b0010001001001011110110111;
      square_table[1909] = 25'b0010001001000111011011000;
      square_table[1910] = 25'b0010001001000010111111001;
      square_table[1911] = 25'b0010001000111110100011110;
      square_table[1912] = 25'b0010001000111010001000011;
      square_table[1913] = 25'b0010001000110101101101011;
      square_table[1914] = 25'b0010001000110001010010100;
      square_table[1915] = 25'b0010001000101100110111111;
      square_table[1916] = 25'b0010001000101000011101011;
      square_table[1917] = 25'b0010001000100100000011001;
      square_table[1918] = 25'b0010001000011111101001010;
      square_table[1919] = 25'b0010001000011011001111100;
      square_table[1920] = 25'b0010001000010110110101110;
      square_table[1921] = 25'b0010001000010010011100011;
      square_table[1922] = 25'b0010001000001110000011010;
      square_table[1923] = 25'b0010001000001001101010011;
      square_table[1924] = 25'b0010001000000101010001101;
      square_table[1925] = 25'b0010001000000000111001000;
      square_table[1926] = 25'b0010000111111100100000110;
      square_table[1927] = 25'b0010000111111000001000101;
      square_table[1928] = 25'b0010000111110011110000111;
      square_table[1929] = 25'b0010000111101111011001001;
      square_table[1930] = 25'b0010000111101011000001101;
      square_table[1931] = 25'b0010000111100110101010011;
      square_table[1932] = 25'b0010000111100010010011011;
      square_table[1933] = 25'b0010000111011101111100101;
      square_table[1934] = 25'b0010000111011001100110000;
      square_table[1935] = 25'b0010000111010101001111100;
      square_table[1936] = 25'b0010000111010000111001010;
      square_table[1937] = 25'b0010000111001100100011010;
      square_table[1938] = 25'b0010000111001000001101100;
      square_table[1939] = 25'b0010000111000011110111111;
      square_table[1940] = 25'b0010000110111111100010101;
      square_table[1941] = 25'b0010000110111011001101100;
      square_table[1942] = 25'b0010000110110110111000011;
      square_table[1943] = 25'b0010000110110010100011110;
      square_table[1944] = 25'b0010000110101110001111001;
      square_table[1945] = 25'b0010000110101001111010111;
      square_table[1946] = 25'b0010000110100101100110110;
      square_table[1947] = 25'b0010000110100001010010110;
      square_table[1948] = 25'b0010000110011100111111001;
      square_table[1949] = 25'b0010000110011000101011101;
      square_table[1950] = 25'b0010000110010100011000011;
      square_table[1951] = 25'b0010000110010000000101001;
      square_table[1952] = 25'b0010000110001011110010011;
      square_table[1953] = 25'b0010000110000111011111110;
      square_table[1954] = 25'b0010000110000011001101010;
      square_table[1955] = 25'b0010000101111110111011000;
      square_table[1956] = 25'b0010000101111010101001000;
      square_table[1957] = 25'b0010000101110110010111001;
      square_table[1958] = 25'b0010000101110010000101100;
      square_table[1959] = 25'b0010000101101101110100000;
      square_table[1960] = 25'b0010000101101001100010110;
      square_table[1961] = 25'b0010000101100101010001110;
      square_table[1962] = 25'b0010000101100001000000111;
      square_table[1963] = 25'b0010000101011100110000010;
      square_table[1964] = 25'b0010000101011000011111111;
      square_table[1965] = 25'b0010000101010100001111101;
      square_table[1966] = 25'b0010000101001111111111101;
      square_table[1967] = 25'b0010000101001011101111110;
      square_table[1968] = 25'b0010000101000111100000010;
      square_table[1969] = 25'b0010000101000011010000110;
      square_table[1970] = 25'b0010000100111111000001101;
      square_table[1971] = 25'b0010000100111010110010101;
      square_table[1972] = 25'b0010000100110110100011111;
      square_table[1973] = 25'b0010000100110010010101010;
      square_table[1974] = 25'b0010000100101110000110110;
      square_table[1975] = 25'b0010000100101001111000101;
      square_table[1976] = 25'b0010000100100101101010110;
      square_table[1977] = 25'b0010000100100001011100111;
      square_table[1978] = 25'b0010000100011101001111010;
      square_table[1979] = 25'b0010000100011001000001111;
      square_table[1980] = 25'b0010000100010100110100101;
      square_table[1981] = 25'b0010000100010000100111110;
      square_table[1982] = 25'b0010000100001100011010111;
      square_table[1983] = 25'b0010000100001000001110010;
      square_table[1984] = 25'b0010000100000100000010000;
      square_table[1985] = 25'b0010000011111111110101110;
      square_table[1986] = 25'b0010000011111011101001110;
      square_table[1987] = 25'b0010000011110111011110000;
      square_table[1988] = 25'b0010000011110011010010011;
      square_table[1989] = 25'b0010000011101111000111000;
      square_table[1990] = 25'b0010000011101010111011111;
      square_table[1991] = 25'b0010000011100110110000110;
      square_table[1992] = 25'b0010000011100010100110000;
      square_table[1993] = 25'b0010000011011110011011011;
      square_table[1994] = 25'b0010000011011010010001000;
      square_table[1995] = 25'b0010000011010110000110111;
      square_table[1996] = 25'b0010000011010001111100111;
      square_table[1997] = 25'b0010000011001101110011000;
      square_table[1998] = 25'b0010000011001001101001011;
      square_table[1999] = 25'b0010000011000101100000000;
      square_table[2000] = 25'b0010000011000001010110110;
      square_table[2001] = 25'b0010000010111101001101111;
      square_table[2002] = 25'b0010000010111001000101000;
      square_table[2003] = 25'b0010000010110100111100011;
      square_table[2004] = 25'b0010000010110000110011111;
      square_table[2005] = 25'b0010000010101100101011110;
      square_table[2006] = 25'b0010000010101000100011101;
      square_table[2007] = 25'b0010000010100100011011110;
      square_table[2008] = 25'b0010000010100000010100001;
      square_table[2009] = 25'b0010000010011100001100101;
      square_table[2010] = 25'b0010000010011000000101100;
      square_table[2011] = 25'b0010000010010011111110011;
      square_table[2012] = 25'b0010000010001111110111100;
      square_table[2013] = 25'b0010000010001011110000110;
      square_table[2014] = 25'b0010000010000111101010011;
      square_table[2015] = 25'b0010000010000011100100000;
      square_table[2016] = 25'b0010000001111111011110000;
      square_table[2017] = 25'b0010000001111011011000001;
      square_table[2018] = 25'b0010000001110111010010010;
      square_table[2019] = 25'b0010000001110011001100111;
      square_table[2020] = 25'b0010000001101111000111100;
      square_table[2021] = 25'b0010000001101011000010011;
      square_table[2022] = 25'b0010000001100110111101011;
      square_table[2023] = 25'b0010000001100010111000110;
      square_table[2024] = 25'b0010000001011110110100001;
      square_table[2025] = 25'b0010000001011010101111111;
      square_table[2026] = 25'b0010000001010110101011101;
      square_table[2027] = 25'b0010000001010010100111101;
      square_table[2028] = 25'b0010000001001110100011111;
      square_table[2029] = 25'b0010000001001010100000010;
      square_table[2030] = 25'b0010000001000110011100111;
      square_table[2031] = 25'b0010000001000010011001101;
      square_table[2032] = 25'b0010000000111110010110101;
      square_table[2033] = 25'b0010000000111010010011110;
      square_table[2034] = 25'b0010000000110110010001001;
      square_table[2035] = 25'b0010000000110010001110101;
      square_table[2036] = 25'b0010000000101110001100011;
      square_table[2037] = 25'b0010000000101010001010010;
      square_table[2038] = 25'b0010000000100110001000011;
      square_table[2039] = 25'b0010000000100010000110110;
      square_table[2040] = 25'b0010000000011110000101010;
      square_table[2041] = 25'b0010000000011010000011111;
      square_table[2042] = 25'b0010000000010110000010110;
      square_table[2043] = 25'b0010000000010010000001111;
      square_table[2044] = 25'b0010000000001110000001001;
      square_table[2045] = 25'b0010000000001010000000100;
      square_table[2046] = 25'b0010000000000110000000001;
      square_table[2047] = 25'b0010000000000010000000000;  
  end
    
  wire [24:0] manx;
  assign manx = {1'b1, mx, 1'b0};  

  logic [24:0] manx_reg;
  logic [24:0] square_reg;
  logic [24:0] twice_reg;
  
  //same to [49:0], because b[49] is definetly 0
  wire [48:0] b;
  assign b = manx_reg * square_reg;

  wire [24:0] m_inv;
  assign m_inv = twice_reg - b[48:24];  //ここでも切り捨ててるけど大丈夫かな？
  
  //基本的にm_invの最上位bitは0になり、次のbitが1になるはずであり、このとき残り23bitを仮数部とすればよい。
  //基本的にはstate==0なはず
  wire state;
  assign state = m_inv[24] ;
  
  wire [7:0] ey;
  assign ey = state ? (8'd254 - ex) : (8'd253 - ex) ;
  
  wire [22:0] my;
  assign my = state ? m_inv[23:1] : m_inv[22:0];
  
  assign y = {sx, ey,  my};

always @(posedge clk) begin
    manx_reg <= manx;
    square_reg <= square_table[x[22:12]];
    twice_reg  <= twice_table[x[22:12]];
end

endmodule   
   
   
   
   
   
   
   
   
   
   
   
   


